netcdf input {
dimensions:
	x = 50 ;
	y = 4 ;
	z = 20 ;
variables:
	double x(x) ;
		x:_FillValue = NaN ;
	double y(y) ;
		y:_FillValue = NaN ;
	double z(z) ;
		z:_FillValue = NaN ;
	double temp(z, y, x) ;
		temp:_FillValue = NaN ;
	double salt(z, y, x) ;
		salt:_FillValue = NaN ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
data:

 x = 2.5, 7.5, 12.5, 17.5, 22.5, 27.5, 32.5, 37.5, 42.5, 47.5, 52.5, 57.5, 
    62.5, 67.5, 72.5, 77.5, 82.5, 87.5, 92.5, 97.5, 102.5, 107.5, 112.5, 
    117.5, 122.5, 127.5, 132.5, 137.5, 142.5, 147.5, 152.5, 157.5, 162.5, 
    167.5, 172.5, 177.5, 182.5, 187.5, 192.5, 197.5, 202.5, 207.5, 212.5, 
    217.5, 222.5, 227.5, 232.5, 237.5, 242.5, 247.5 ;

 y = 2.5, 7.5, 12.5, 17.5 ;

 z = 12.5, 37.5, 62.5, 87.5, 112.5, 137.5, 162.5, 187.5, 212.5, 237.5, 262.5, 
    287.5, 312.5, 337.5, 362.5, 387.5, 412.5, 437.5, 462.5, 487.5 ;

 temp =
  19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8190423302543, 
    19.7705519423679, 19.7238599875462, 19.6801161766785, 19.6403976275658, 
    19.6056823427057, 19.5768251276247, 19.5545365427297, 19.5393654069525, 
    19.531685284006, 19.531685284006, 19.5393654069525, 19.5545365427297, 
    19.5768251276247, 19.6056823427057, 19.6403976275658, 19.6801161766785, 
    19.7238599875462, 19.7705519423679, 19.8190423302543, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897,
  19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8190423302543, 
    19.7705519423679, 19.7238599875462, 19.6801161766785, 19.6403976275658, 
    19.6056823427057, 19.5768251276247, 19.5545365427297, 19.5393654069525, 
    19.531685284006, 19.531685284006, 19.5393654069525, 19.5545365427297, 
    19.5768251276247, 19.6056823427057, 19.6403976275658, 19.6801161766785, 
    19.7238599875462, 19.7705519423679, 19.8190423302543, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897,
  19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8190423302543, 
    19.7705519423679, 19.7238599875462, 19.6801161766785, 19.6403976275658, 
    19.6056823427057, 19.5768251276247, 19.5545365427297, 19.5393654069525, 
    19.531685284006, 19.531685284006, 19.5393654069525, 19.5545365427297, 
    19.5768251276247, 19.6056823427057, 19.6403976275658, 19.6801161766785, 
    19.7238599875462, 19.7705519423679, 19.8190423302543, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897,
  19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8190423302543, 
    19.7705519423679, 19.7238599875462, 19.6801161766785, 19.6403976275658, 
    19.6056823427057, 19.5768251276247, 19.5545365427297, 19.5393654069525, 
    19.531685284006, 19.531685284006, 19.5393654069525, 19.5545365427297, 
    19.5768251276247, 19.6056823427057, 19.6403976275658, 19.6801161766785, 
    19.7238599875462, 19.7705519423679, 19.8190423302543, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897,
  19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.2822788428828, 
    19.1864920613902, 19.0942578626361, 19.0078473587017, 18.9293882629739, 
    18.8608124987802, 18.8038086290251, 18.7597802781669, 18.7298115703254, 
    18.7146404345482, 18.7146404345482, 18.7298115703254, 18.7597802781669, 
    18.8038086290251, 18.8608124987802, 18.9293882629739, 19.0078473587017, 
    19.0942578626361, 19.1864920613902, 19.2822788428828, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692,
  19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.2822788428828, 
    19.1864920613902, 19.0942578626361, 19.0078473587017, 18.9293882629739, 
    18.8608124987802, 18.8038086290251, 18.7597802781669, 18.7298115703254, 
    18.7146404345482, 18.7146404345482, 18.7298115703254, 18.7597802781669, 
    18.8038086290251, 18.8608124987802, 18.9293882629739, 19.0078473587017, 
    19.0942578626361, 19.1864920613902, 19.2822788428828, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692,
  19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.2822788428828, 
    19.1864920613902, 19.0942578626361, 19.0078473587017, 18.9293882629739, 
    18.8608124987802, 18.8038086290251, 18.7597802781669, 18.7298115703254, 
    18.7146404345482, 18.7146404345482, 18.7298115703254, 18.7597802781669, 
    18.8038086290251, 18.8608124987802, 18.9293882629739, 19.0078473587017, 
    19.0942578626361, 19.1864920613902, 19.2822788428828, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692,
  19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.2822788428828, 
    19.1864920613902, 19.0942578626361, 19.0078473587017, 18.9293882629739, 
    18.8608124987802, 18.8038086290251, 18.7597802781669, 18.7298115703254, 
    18.7146404345482, 18.7146404345482, 18.7298115703254, 18.7597802781669, 
    18.8038086290251, 18.8608124987802, 18.9293882629739, 19.0078473587017, 
    19.0942578626361, 19.1864920613902, 19.2822788428828, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692,
  18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.7467093497915, 
    18.6059847631511, 18.4704794325458, 18.3435299489315, 18.2282622299161, 
    18.1275145492933, 18.0437676493225, 17.9790836566208, 17.9350553057626, 
    17.9127667208677, 17.9127667208677, 17.9350553057626, 17.9790836566208, 
    18.0437676493225, 18.1275145492933, 18.2282622299161, 18.3435299489315, 
    18.4704794325458, 18.6059847631511, 18.7467093497915, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487,
  18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.7467093497915, 
    18.6059847631511, 18.4704794325458, 18.3435299489315, 18.2282622299161, 
    18.1275145492933, 18.0437676493225, 17.9790836566208, 17.9350553057626, 
    17.9127667208677, 17.9127667208677, 17.9350553057626, 17.9790836566208, 
    18.0437676493225, 18.1275145492933, 18.2282622299161, 18.3435299489315, 
    18.4704794325458, 18.6059847631511, 18.7467093497915, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487,
  18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.7467093497915, 
    18.6059847631511, 18.4704794325458, 18.3435299489315, 18.2282622299161, 
    18.1275145492933, 18.0437676493225, 17.9790836566208, 17.9350553057626, 
    17.9127667208677, 17.9127667208677, 17.9350553057626, 17.9790836566208, 
    18.0437676493225, 18.1275145492933, 18.2282622299161, 18.3435299489315, 
    18.4704794325458, 18.6059847631511, 18.7467093497915, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487,
  18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.7467093497915, 
    18.6059847631511, 18.4704794325458, 18.3435299489315, 18.2282622299161, 
    18.1275145492933, 18.0437676493225, 17.9790836566208, 17.9350553057626, 
    17.9127667208677, 17.9127667208677, 17.9350553057626, 17.9790836566208, 
    18.0437676493225, 18.1275145492933, 18.2282622299161, 18.3435299489315, 
    18.4704794325458, 18.6059847631511, 18.7467093497915, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487,
  18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.2128940063741, 
    18.0306967209471, 17.8552568494465, 17.6908943037602, 17.541656235251, 
    17.4112173804584, 17.3027895768891, 17.2190426769182, 17.1620388071631, 
    17.1331815920821, 17.1331815920821, 17.1620388071631, 17.2190426769182, 
    17.3027895768891, 17.4112173804584, 17.541656235251, 17.6908943037602, 
    17.8552568494465, 18.0306967209471, 18.2128940063741, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282,
  18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.2128940063741, 
    18.0306967209471, 17.8552568494465, 17.6908943037602, 17.541656235251, 
    17.4112173804584, 17.3027895768891, 17.2190426769182, 17.1620388071631, 
    17.1331815920821, 17.1331815920821, 17.1620388071631, 17.2190426769182, 
    17.3027895768891, 17.4112173804584, 17.541656235251, 17.6908943037602, 
    17.8552568494465, 18.0306967209471, 18.2128940063741, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282,
  18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.2128940063741, 
    18.0306967209471, 17.8552568494465, 17.6908943037602, 17.541656235251, 
    17.4112173804584, 17.3027895768891, 17.2190426769182, 17.1620388071631, 
    17.1331815920821, 17.1331815920821, 17.1620388071631, 17.2190426769182, 
    17.3027895768891, 17.4112173804584, 17.541656235251, 17.6908943037602, 
    17.8552568494465, 18.0306967209471, 18.2128940063741, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282,
  18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.2128940063741, 
    18.0306967209471, 17.8552568494465, 17.6908943037602, 17.541656235251, 
    17.4112173804584, 17.3027895768891, 17.2190426769182, 17.1620388071631, 
    17.1331815920821, 17.1331815920821, 17.1620388071631, 17.2190426769182, 
    17.3027895768891, 17.4112173804584, 17.541656235251, 17.6908943037602, 
    17.8552568494465, 18.0306967209471, 18.2128940063741, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282,
  17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.6813497750378, 
    17.4621660926696, 17.2511115921615, 17.0533831357659, 16.8738494543024, 
    16.7169312628467, 16.5864924080541, 16.4857447274313, 16.4171689632377, 
    16.3824536783775, 16.3824536783775, 16.4171689632377, 16.4857447274313, 
    16.5864924080541, 16.7169312628467, 16.8738494543024, 17.0533831357659, 
    17.2511115921615, 17.4621660926696, 17.6813497750378, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077,
  17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.6813497750378, 
    17.4621660926696, 17.2511115921615, 17.0533831357659, 16.8738494543024, 
    16.7169312628467, 16.5864924080541, 16.4857447274313, 16.4171689632377, 
    16.3824536783775, 16.3824536783775, 16.4171689632377, 16.4857447274313, 
    16.5864924080541, 16.7169312628467, 16.8738494543024, 17.0533831357659, 
    17.2511115921615, 17.4621660926696, 17.6813497750378, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077,
  17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.6813497750378, 
    17.4621660926696, 17.2511115921615, 17.0533831357659, 16.8738494543024, 
    16.7169312628467, 16.5864924080541, 16.4857447274313, 16.4171689632377, 
    16.3824536783775, 16.3824536783775, 16.4171689632377, 16.4857447274313, 
    16.5864924080541, 16.7169312628467, 16.8738494543024, 17.0533831357659, 
    17.2511115921615, 17.4621660926696, 17.6813497750378, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077,
  17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.6813497750378, 
    17.4621660926696, 17.2511115921615, 17.0533831357659, 16.8738494543024, 
    16.7169312628467, 16.5864924080541, 16.4857447274313, 16.4171689632377, 
    16.3824536783775, 16.3824536783775, 16.4171689632377, 16.4857447274313, 
    16.5864924080541, 16.7169312628467, 16.8738494543024, 17.0533831357659, 
    17.2511115921615, 17.4621660926696, 17.6813497750378, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077,
  17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.1525376958729, 
    16.9017646462522, 16.660292378989, 16.4340667427037, 16.2286581633617, 
    16.0491244818981, 15.899886413389, 15.7846186943736, 15.7061595986457, 
    15.6664410495331, 15.6664410495331, 15.7061595986457, 15.7846186943736, 
    15.899886413389, 16.0491244818981, 16.2286581633617, 16.4340667427037, 
    16.660292378989, 16.9017646462522, 17.1525376958729, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872,
  17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.1525376958729, 
    16.9017646462522, 16.660292378989, 16.4340667427037, 16.2286581633617, 
    16.0491244818981, 15.899886413389, 15.7846186943736, 15.7061595986457, 
    15.6664410495331, 15.6664410495331, 15.7061595986457, 15.7846186943736, 
    15.899886413389, 16.0491244818981, 16.2286581633617, 16.4340667427037, 
    16.660292378989, 16.9017646462522, 17.1525376958729, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872,
  17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.1525376958729, 
    16.9017646462522, 16.660292378989, 16.4340667427037, 16.2286581633617, 
    16.0491244818981, 15.899886413389, 15.7846186943736, 15.7061595986457, 
    15.6664410495331, 15.6664410495331, 15.7061595986457, 15.7846186943736, 
    15.899886413389, 16.0491244818981, 16.2286581633617, 16.4340667427037, 
    16.660292378989, 16.9017646462522, 17.1525376958729, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872,
  17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.1525376958729, 
    16.9017646462522, 16.660292378989, 16.4340667427037, 16.2286581633617, 
    16.0491244818981, 15.899886413389, 15.7846186943736, 15.7061595986457, 
    15.6664410495331, 15.6664410495331, 15.7061595986457, 15.7846186943736, 
    15.899886413389, 16.0491244818981, 16.2286581633617, 16.4340667427037, 
    16.660292378989, 16.9017646462522, 17.1525376958729, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872,
  16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.6268515343158, 
    16.3506639821924, 16.0847197967945, 15.8355674065847, 15.6093417702995, 
    15.4116133139039, 15.2472507682176, 15.1203012846034, 15.033890780669, 
    14.9901469698013, 14.9901469698013, 15.033890780669, 15.1203012846034, 
    15.2472507682176, 15.4116133139039, 15.6093417702995, 15.8355674065847, 
    16.0847197967945, 16.3506639821924, 16.6268515343158, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667,
  16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.6268515343158, 
    16.3506639821924, 16.0847197967945, 15.8355674065847, 15.6093417702995, 
    15.4116133139039, 15.2472507682176, 15.1203012846034, 15.033890780669, 
    14.9901469698013, 14.9901469698013, 15.033890780669, 15.1203012846034, 
    15.2472507682176, 15.4116133139039, 15.6093417702995, 15.8355674065847, 
    16.0847197967945, 16.3506639821924, 16.6268515343158, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667,
  16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.6268515343158, 
    16.3506639821924, 16.0847197967945, 15.8355674065847, 15.6093417702995, 
    15.4116133139039, 15.2472507682176, 15.1203012846034, 15.033890780669, 
    14.9901469698013, 14.9901469698013, 15.033890780669, 15.1203012846034, 
    15.2472507682176, 15.4116133139039, 15.6093417702995, 15.8355674065847, 
    16.0847197967945, 16.3506639821924, 16.6268515343158, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667,
  16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.6268515343158, 
    16.3506639821924, 16.0847197967945, 15.8355674065847, 15.6093417702995, 
    15.4116133139039, 15.2472507682176, 15.1203012846034, 15.033890780669, 
    14.9901469698013, 14.9901469698013, 15.033890780669, 15.1203012846034, 
    15.2472507682176, 15.4116133139039, 15.6093417702995, 15.8355674065847, 
    16.0847197967945, 16.3506639821924, 16.6268515343158, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667,
  16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.104608085337, 
    15.8098066848581, 15.5259390097881, 15.2599948243902, 15.018522557127, 
    14.8074680566189, 14.6320281851183, 14.496522854513, 14.4042886557589, 
    14.3575967009372, 14.3575967009372, 14.4042886557589, 14.496522854513, 
    14.6320281851183, 14.8074680566189, 15.018522557127, 15.2599948243902, 
    15.5259390097881, 15.8098066848581, 16.104608085337, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462,
  16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.104608085337, 
    15.8098066848581, 15.5259390097881, 15.2599948243902, 15.018522557127, 
    14.8074680566189, 14.6320281851183, 14.496522854513, 14.4042886557589, 
    14.3575967009372, 14.3575967009372, 14.4042886557589, 14.496522854513, 
    14.6320281851183, 14.8074680566189, 15.018522557127, 15.2599948243902, 
    15.5259390097881, 15.8098066848581, 16.104608085337, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462,
  16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.104608085337, 
    15.8098066848581, 15.5259390097881, 15.2599948243902, 15.018522557127, 
    14.8074680566189, 14.6320281851183, 14.496522854513, 14.4042886557589, 
    14.3575967009372, 14.3575967009372, 14.4042886557589, 14.496522854513, 
    14.6320281851183, 14.8074680566189, 15.018522557127, 15.2599948243902, 
    15.5259390097881, 15.8098066848581, 16.104608085337, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462,
  16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.104608085337, 
    15.8098066848581, 15.5259390097881, 15.2599948243902, 15.018522557127, 
    14.8074680566189, 14.6320281851183, 14.496522854513, 14.4042886557589, 
    14.3575967009372, 14.3575967009372, 14.4042886557589, 14.496522854513, 
    14.6320281851183, 14.8074680566189, 15.018522557127, 15.2599948243902, 
    15.5259390097881, 15.8098066848581, 16.104608085337, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462,
  15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.5860393728976, 
    15.2798831129327, 14.9850817124538, 14.7088941603304, 14.4581211107097, 
    14.2389374283414, 14.0567401429143, 13.9160155562739, 13.8202287747812, 
    13.7717383868948, 13.7717383868948, 13.8202287747812, 13.9160155562739, 
    14.0567401429143, 14.2389374283414, 14.4581211107097, 14.7088941603304, 
    14.9850817124538, 15.2798831129327, 15.5860393728976, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256,
  15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.5860393728976, 
    15.2798831129327, 14.9850817124538, 14.7088941603304, 14.4581211107097, 
    14.2389374283414, 14.0567401429143, 13.9160155562739, 13.8202287747812, 
    13.7717383868948, 13.7717383868948, 13.8202287747812, 13.9160155562739, 
    14.0567401429143, 14.2389374283414, 14.4581211107097, 14.7088941603304, 
    14.9850817124538, 15.2798831129327, 15.5860393728976, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256,
  15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.5860393728976, 
    15.2798831129327, 14.9850817124538, 14.7088941603304, 14.4581211107097, 
    14.2389374283414, 14.0567401429143, 13.9160155562739, 13.8202287747812, 
    13.7717383868948, 13.7717383868948, 13.8202287747812, 13.9160155562739, 
    14.0567401429143, 14.2389374283414, 14.4581211107097, 14.7088941603304, 
    14.9850817124538, 15.2798831129327, 15.5860393728976, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256,
  15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.5860393728976, 
    15.2798831129327, 14.9850817124538, 14.7088941603304, 14.4581211107097, 
    14.2389374283414, 14.0567401429143, 13.9160155562739, 13.8202287747812, 
    13.7717383868948, 13.7717383868948, 13.8202287747812, 13.9160155562739, 
    14.0567401429143, 14.2389374283414, 14.4581211107097, 14.7088941603304, 
    14.9850817124538, 15.2798831129327, 15.5860393728976, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256,
  15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.0712869367494, 
    14.7613144004933, 14.4628382634749, 14.1832079987732, 13.9293090315448, 
    13.7073931970051, 13.5229247994969, 13.3804460631826, 13.2834652874098, 
    13.2343704607389, 13.2343704607389, 13.2834652874098, 13.3804460631826, 
    13.5229247994969, 13.7073931970051, 13.9293090315448, 14.1832079987732, 
    14.4628382634749, 14.7613144004933, 15.0712869367494, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051,
  15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.0712869367494, 
    14.7613144004933, 14.4628382634749, 14.1832079987732, 13.9293090315448, 
    13.7073931970051, 13.5229247994969, 13.3804460631826, 13.2834652874098, 
    13.2343704607389, 13.2343704607389, 13.2834652874098, 13.3804460631826, 
    13.5229247994969, 13.7073931970051, 13.9293090315448, 14.1832079987732, 
    14.4628382634749, 14.7613144004933, 15.0712869367494, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051,
  15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.0712869367494, 
    14.7613144004933, 14.4628382634749, 14.1832079987732, 13.9293090315448, 
    13.7073931970051, 13.5229247994969, 13.3804460631826, 13.2834652874098, 
    13.2343704607389, 13.2343704607389, 13.2834652874098, 13.3804460631826, 
    13.5229247994969, 13.7073931970051, 13.9293090315448, 14.1832079987732, 
    14.4628382634749, 14.7613144004933, 15.0712869367494, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051,
  15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.0712869367494, 
    14.7613144004933, 14.4628382634749, 14.1832079987732, 13.9293090315448, 
    13.7073931970051, 13.5229247994969, 13.3804460631826, 13.2834652874098, 
    13.2343704607389, 13.2343704607389, 13.2834652874098, 13.3804460631826, 
    13.5229247994969, 13.7073931970051, 13.9293090315448, 14.1832079987732, 
    14.4628382634749, 14.7613144004933, 15.0712869367494, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051,
  14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.5603983472566, 
    14.2542420872917, 13.9594406868128, 13.6832531346893, 13.4324800850686, 
    13.2132964027003, 13.0310991172733, 12.8903745306328, 12.7945877491402, 
    12.7460973612538, 12.7460973612538, 12.7945877491402, 12.8903745306328, 
    13.0310991172733, 13.2132964027003, 13.4324800850686, 13.6832531346893, 
    13.9594406868128, 14.2542420872917, 14.5603983472566, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846,
  14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.5603983472566, 
    14.2542420872917, 13.9594406868128, 13.6832531346893, 13.4324800850686, 
    13.2132964027003, 13.0310991172733, 12.8903745306328, 12.7945877491402, 
    12.7460973612538, 12.7460973612538, 12.7945877491402, 12.8903745306328, 
    13.0310991172733, 13.2132964027003, 13.4324800850686, 13.6832531346893, 
    13.9594406868128, 14.2542420872917, 14.5603983472566, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846,
  14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.5603983472566, 
    14.2542420872917, 13.9594406868128, 13.6832531346893, 13.4324800850686, 
    13.2132964027003, 13.0310991172733, 12.8903745306328, 12.7945877491402, 
    12.7460973612538, 12.7460973612538, 12.7945877491402, 12.8903745306328, 
    13.0310991172733, 13.2132964027003, 13.4324800850686, 13.6832531346893, 
    13.9594406868128, 14.2542420872917, 14.5603983472566, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846,
  14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.5603983472566, 
    14.2542420872917, 13.9594406868128, 13.6832531346893, 13.4324800850686, 
    13.2132964027003, 13.0310991172733, 12.8903745306328, 12.7945877491402, 
    12.7460973612538, 12.7460973612538, 12.7945877491402, 12.8903745306328, 
    13.0310991172733, 13.2132964027003, 13.4324800850686, 13.6832531346893, 
    13.9594406868128, 14.2542420872917, 14.5603983472566, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846,
  14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.0533260340549, 
    13.758524633576, 13.4746569585061, 13.2087127731082, 12.9672405058449, 
    12.7561860053369, 12.5807461338362, 12.4452408032309, 12.3530066044769, 
    12.3063146496551, 12.3063146496551, 12.3530066044769, 12.4452408032309, 
    12.5807461338362, 12.7561860053369, 12.9672405058449, 13.2087127731082, 
    13.4746569585061, 13.758524633576, 14.0533260340549, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641,
  14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.0533260340549, 
    13.758524633576, 13.4746569585061, 13.2087127731082, 12.9672405058449, 
    12.7561860053369, 12.5807461338362, 12.4452408032309, 12.3530066044769, 
    12.3063146496551, 12.3063146496551, 12.3530066044769, 12.4452408032309, 
    12.5807461338362, 12.7561860053369, 12.9672405058449, 13.2087127731082, 
    13.4746569585061, 13.758524633576, 14.0533260340549, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641,
  14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.0533260340549, 
    13.758524633576, 13.4746569585061, 13.2087127731082, 12.9672405058449, 
    12.7561860053369, 12.5807461338362, 12.4452408032309, 12.3530066044769, 
    12.3063146496551, 12.3063146496551, 12.3530066044769, 12.4452408032309, 
    12.5807461338362, 12.7561860053369, 12.9672405058449, 13.2087127731082, 
    13.4746569585061, 13.758524633576, 14.0533260340549, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641,
  14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.0533260340549, 
    13.758524633576, 13.4746569585061, 13.2087127731082, 12.9672405058449, 
    12.7561860053369, 12.5807461338362, 12.4452408032309, 12.3530066044769, 
    12.3063146496551, 12.3063146496551, 12.3530066044769, 12.4452408032309, 
    12.5807461338362, 12.7561860053369, 12.9672405058449, 13.2087127731082, 
    13.4746569585061, 13.758524633576, 14.0533260340549, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641,
  13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.5499284573927, 
    13.2737409052693, 13.0077967198714, 12.7586443296617, 12.5324186933764, 
    12.3346902369808, 12.1703276912945, 12.0433782076803, 11.9569677037459, 
    11.9132238928782, 11.9132238928782, 11.9569677037459, 12.0433782076803, 
    12.1703276912945, 12.3346902369808, 12.5324186933764, 12.7586443296617, 
    13.0077967198714, 13.2737409052693, 13.5499284573927, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436,
  13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.5499284573927, 
    13.2737409052693, 13.0077967198714, 12.7586443296617, 12.5324186933764, 
    12.3346902369808, 12.1703276912945, 12.0433782076803, 11.9569677037459, 
    11.9132238928782, 11.9132238928782, 11.9569677037459, 12.0433782076803, 
    12.1703276912945, 12.3346902369808, 12.5324186933764, 12.7586443296617, 
    13.0077967198714, 13.2737409052693, 13.5499284573927, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436,
  13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.5499284573927, 
    13.2737409052693, 13.0077967198714, 12.7586443296617, 12.5324186933764, 
    12.3346902369808, 12.1703276912945, 12.0433782076803, 11.9569677037459, 
    11.9132238928782, 11.9132238928782, 11.9569677037459, 12.0433782076803, 
    12.1703276912945, 12.3346902369808, 12.5324186933764, 12.7586443296617, 
    13.0077967198714, 13.2737409052693, 13.5499284573927, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436,
  13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.5499284573927, 
    13.2737409052693, 13.0077967198714, 12.7586443296617, 12.5324186933764, 
    12.3346902369808, 12.1703276912945, 12.0433782076803, 11.9569677037459, 
    11.9132238928782, 11.9132238928782, 11.9569677037459, 12.0433782076803, 
    12.1703276912945, 12.3346902369808, 12.5324186933764, 12.7586443296617, 
    13.0077967198714, 13.2737409052693, 13.5499284573927, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436,
  13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.0499735933088, 
    12.7992005436881, 12.5577282764249, 12.3315026401396, 12.1260940607976, 
    11.946560379334, 11.7973223108249, 11.6820545918095, 11.6035954960816, 
    11.563876946969, 11.563876946969, 11.6035954960816, 11.6820545918095, 
    11.7973223108249, 11.946560379334, 12.1260940607976, 12.3315026401396, 
    12.5577282764249, 12.7992005436881, 13.0499735933088, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231,
  13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.0499735933088, 
    12.7992005436881, 12.5577282764249, 12.3315026401396, 12.1260940607976, 
    11.946560379334, 11.7973223108249, 11.6820545918095, 11.6035954960816, 
    11.563876946969, 11.563876946969, 11.6035954960816, 11.6820545918095, 
    11.7973223108249, 11.946560379334, 12.1260940607976, 12.3315026401396, 
    12.5577282764249, 12.7992005436881, 13.0499735933088, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231,
  13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.0499735933088, 
    12.7992005436881, 12.5577282764249, 12.3315026401396, 12.1260940607976, 
    11.946560379334, 11.7973223108249, 11.6820545918095, 11.6035954960816, 
    11.563876946969, 11.563876946969, 11.6035954960816, 11.6820545918095, 
    11.7973223108249, 11.946560379334, 12.1260940607976, 12.3315026401396, 
    12.5577282764249, 12.7992005436881, 13.0499735933088, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231,
  13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.0499735933088, 
    12.7992005436881, 12.5577282764249, 12.3315026401396, 12.1260940607976, 
    11.946560379334, 11.7973223108249, 11.6820545918095, 11.6035954960816, 
    11.563876946969, 11.563876946969, 11.6035954960816, 11.6820545918095, 
    11.7973223108249, 11.946560379334, 12.1260940607976, 12.3315026401396, 
    12.5577282764249, 12.7992005436881, 13.0499735933088, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231,
  12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.5531446468327, 
    12.3339609644644, 12.1229064639564, 11.9251780075608, 11.7456443260973, 
    11.5887261346416, 11.458287279849, 11.3575395992262, 11.2889638350325, 
    11.2542485501723, 11.2542485501723, 11.2889638350325, 11.3575395992262, 
    11.458287279849, 11.5887261346416, 11.7456443260973, 11.9251780075608, 
    12.1229064639564, 12.3339609644644, 12.5531446468327, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026,
  12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.5531446468327, 
    12.3339609644644, 12.1229064639564, 11.9251780075608, 11.7456443260973, 
    11.5887261346416, 11.458287279849, 11.3575395992262, 11.2889638350325, 
    11.2542485501723, 11.2542485501723, 11.2889638350325, 11.3575395992262, 
    11.458287279849, 11.5887261346416, 11.7456443260973, 11.9251780075608, 
    12.1229064639564, 12.3339609644644, 12.5531446468327, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026,
  12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.5531446468327, 
    12.3339609644644, 12.1229064639564, 11.9251780075608, 11.7456443260973, 
    11.5887261346416, 11.458287279849, 11.3575395992262, 11.2889638350325, 
    11.2542485501723, 11.2542485501723, 11.2889638350325, 11.3575395992262, 
    11.458287279849, 11.5887261346416, 11.7456443260973, 11.9251780075608, 
    12.1229064639564, 12.3339609644644, 12.5531446468327, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026,
  12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.5531446468327, 
    12.3339609644644, 12.1229064639564, 11.9251780075608, 11.7456443260973, 
    11.5887261346416, 11.458287279849, 11.3575395992262, 11.2889638350325, 
    11.2542485501723, 11.2542485501723, 11.2889638350325, 11.3575395992262, 
    11.458287279849, 11.5887261346416, 11.7456443260973, 11.9251780075608, 
    12.1229064639564, 12.3339609644644, 12.5531446468327, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026,
  12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.059047852528, 
    11.8768505671009, 11.7014106956003, 11.537048149914, 11.3878100814048, 
    11.2573712266122, 11.1489434230429, 11.0651965230721, 11.0081926533169, 
    10.9793354382359, 10.9793354382359, 11.0081926533169, 11.0651965230721, 
    11.1489434230429, 11.2573712266122, 11.3878100814048, 11.537048149914, 
    11.7014106956003, 11.8768505671009, 12.059047852528, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821,
  12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.059047852528, 
    11.8768505671009, 11.7014106956003, 11.537048149914, 11.3878100814048, 
    11.2573712266122, 11.1489434230429, 11.0651965230721, 11.0081926533169, 
    10.9793354382359, 10.9793354382359, 11.0081926533169, 11.0651965230721, 
    11.1489434230429, 11.2573712266122, 11.3878100814048, 11.537048149914, 
    11.7014106956003, 11.8768505671009, 12.059047852528, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821,
  12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.059047852528, 
    11.8768505671009, 11.7014106956003, 11.537048149914, 11.3878100814048, 
    11.2573712266122, 11.1489434230429, 11.0651965230721, 11.0081926533169, 
    10.9793354382359, 10.9793354382359, 11.0081926533169, 11.0651965230721, 
    11.1489434230429, 11.2573712266122, 11.3878100814048, 11.537048149914, 
    11.7014106956003, 11.8768505671009, 12.059047852528, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821,
  12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.059047852528, 
    11.8768505671009, 11.7014106956003, 11.537048149914, 11.3878100814048, 
    11.2573712266122, 11.1489434230429, 11.0651965230721, 11.0081926533169, 
    10.9793354382359, 10.9793354382359, 11.0081926533169, 11.0651965230721, 
    11.1489434230429, 11.2573712266122, 11.3878100814048, 11.537048149914, 
    11.7014106956003, 11.8768505671009, 12.059047852528, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821,
  11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.5672221703043, 
    11.4264975836639, 11.2909922530586, 11.1640427694444, 11.048775050429, 
    10.9480273698062, 10.8642804698353, 10.7995964771337, 10.7555681262754, 
    10.7332795413805, 10.7332795413805, 10.7555681262754, 10.7995964771337, 
    10.8642804698353, 10.9480273698062, 11.048775050429, 11.1640427694444, 
    11.2909922530586, 11.4264975836639, 11.5672221703043, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615,
  11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.5672221703043, 
    11.4264975836639, 11.2909922530586, 11.1640427694444, 11.048775050429, 
    10.9480273698062, 10.8642804698353, 10.7995964771337, 10.7555681262754, 
    10.7332795413805, 10.7332795413805, 10.7555681262754, 10.7995964771337, 
    10.8642804698353, 10.9480273698062, 11.048775050429, 11.1640427694444, 
    11.2909922530586, 11.4264975836639, 11.5672221703043, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615,
  11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.5672221703043, 
    11.4264975836639, 11.2909922530586, 11.1640427694444, 11.048775050429, 
    10.9480273698062, 10.8642804698353, 10.7995964771337, 10.7555681262754, 
    10.7332795413805, 10.7332795413805, 10.7555681262754, 10.7995964771337, 
    10.8642804698353, 10.9480273698062, 11.048775050429, 11.1640427694444, 
    11.2909922530586, 11.4264975836639, 11.5672221703043, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615,
  11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.5672221703043, 
    11.4264975836639, 11.2909922530586, 11.1640427694444, 11.048775050429, 
    10.9480273698062, 10.8642804698353, 10.7995964771337, 10.7555681262754, 
    10.7332795413805, 10.7332795413805, 10.7555681262754, 10.7995964771337, 
    10.8642804698353, 10.9480273698062, 11.048775050429, 11.1640427694444, 
    11.2909922530586, 11.4264975836639, 11.5672221703043, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615,
  11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.0771506377546, 
    10.981363856262, 10.8891296575079, 10.8027191535735, 10.7242600578457, 
    10.655684293652, 10.5986804238969, 10.5546520730387, 10.5246833651972, 
    10.50951222942, 10.50951222942, 10.5246833651972, 10.5546520730387, 
    10.5986804238969, 10.655684293652, 10.7242600578457, 10.8027191535735, 
    10.8891296575079, 10.981363856262, 11.0771506377546, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641,
  11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.0771506377546, 
    10.981363856262, 10.8891296575079, 10.8027191535735, 10.7242600578457, 
    10.655684293652, 10.5986804238969, 10.5546520730387, 10.5246833651972, 
    10.50951222942, 10.50951222942, 10.5246833651972, 10.5546520730387, 
    10.5986804238969, 10.655684293652, 10.7242600578457, 10.8027191535735, 
    10.8891296575079, 10.981363856262, 11.0771506377546, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641,
  11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.0771506377546, 
    10.981363856262, 10.8891296575079, 10.8027191535735, 10.7242600578457, 
    10.655684293652, 10.5986804238969, 10.5546520730387, 10.5246833651972, 
    10.50951222942, 10.50951222942, 10.5246833651972, 10.5546520730387, 
    10.5986804238969, 10.655684293652, 10.7242600578457, 10.8027191535735, 
    10.8891296575079, 10.981363856262, 11.0771506377546, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641,
  11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.0771506377546, 
    10.981363856262, 10.8891296575079, 10.8027191535735, 10.7242600578457, 
    10.655684293652, 10.5986804238969, 10.5546520730387, 10.5246833651972, 
    10.50951222942, 10.50951222942, 10.5246833651972, 10.5546520730387, 
    10.5986804238969, 10.655684293652, 10.7242600578457, 10.8027191535735, 
    10.8891296575079, 10.981363856262, 11.0771506377546, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641,
  10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.5882730994851, 
    10.5397827115987, 10.4930907567769, 10.4493469459093, 10.4096283967966, 
    10.3749131119364, 10.3460558968554, 10.3237673119605, 10.3085961761833, 
    10.3009160532368, 10.3009160532368, 10.3085961761833, 10.3237673119605, 
    10.3460558968554, 10.3749131119364, 10.4096283967966, 10.4493469459093, 
    10.4930907567769, 10.5397827115987, 10.5882730994851, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205,
  10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.5882730994851, 
    10.5397827115987, 10.4930907567769, 10.4493469459093, 10.4096283967966, 
    10.3749131119364, 10.3460558968554, 10.3237673119605, 10.3085961761833, 
    10.3009160532368, 10.3009160532368, 10.3085961761833, 10.3237673119605, 
    10.3460558968554, 10.3749131119364, 10.4096283967966, 10.4493469459093, 
    10.4930907567769, 10.5397827115987, 10.5882730994851, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205,
  10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.5882730994851, 
    10.5397827115987, 10.4930907567769, 10.4493469459093, 10.4096283967966, 
    10.3749131119364, 10.3460558968554, 10.3237673119605, 10.3085961761833, 
    10.3009160532368, 10.3009160532368, 10.3085961761833, 10.3237673119605, 
    10.3460558968554, 10.3749131119364, 10.4096283967966, 10.4493469459093, 
    10.4930907567769, 10.5397827115987, 10.5882730994851, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205,
  10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.5882730994851, 
    10.5397827115987, 10.4930907567769, 10.4493469459093, 10.4096283967966, 
    10.3749131119364, 10.3460558968554, 10.3237673119605, 10.3085961761833, 
    10.3009160532368, 10.3009160532368, 10.3085961761833, 10.3237673119605, 
    10.3460558968554, 10.3749131119364, 10.4096283967966, 10.4493469459093, 
    10.4930907567769, 10.5397827115987, 10.5882730994851, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205,
  10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1,
  10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1,
  10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1,
  10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1 ;

 salt =
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35 ;
}
