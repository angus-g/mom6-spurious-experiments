netcdf input_rho {
dimensions:
	x = 128 ;
	y = 4 ;
	z = 20 ;
variables:
	double x(x) ;
		x:_FillValue = NaN ;
	double y(y) ;
		y:_FillValue = NaN ;
	double z(z) ;
		z:_FillValue = NaN ;
	double temp(z, y, x) ;
		temp:_FillValue = NaN ;
	double salt(z, y, x) ;
		salt:_FillValue = NaN ;
	double h(z, y, x) ;
		h:_FillValue = NaN ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
data:

 x = 250, 750, 1250, 1750, 2250, 2750, 3250, 3750, 4250, 4750, 5250, 5750, 
    6250, 6750, 7250, 7750, 8250, 8750, 9250, 9750, 10250, 10750, 11250, 
    11750, 12250, 12750, 13250, 13750, 14250, 14750, 15250, 15750, 16250, 
    16750, 17250, 17750, 18250, 18750, 19250, 19750, 20250, 20750, 21250, 
    21750, 22250, 22750, 23250, 23750, 24250, 24750, 25250, 25750, 26250, 
    26750, 27250, 27750, 28250, 28750, 29250, 29750, 30250, 30750, 31250, 
    31750, 32250, 32750, 33250, 33750, 34250, 34750, 35250, 35750, 36250, 
    36750, 37250, 37750, 38250, 38750, 39250, 39750, 40250, 40750, 41250, 
    41750, 42250, 42750, 43250, 43750, 44250, 44750, 45250, 45750, 46250, 
    46750, 47250, 47750, 48250, 48750, 49250, 49750, 50250, 50750, 51250, 
    51750, 52250, 52750, 53250, 53750, 54250, 54750, 55250, 55750, 56250, 
    56750, 57250, 57750, 58250, 58750, 59250, 59750, 60250, 60750, 61250, 
    61750, 62250, 62750, 63250, 63750 ;

 y = 0, 1, 2, 3 ;

 z = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19 ;

 temp =
  30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30,
  30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30,
  30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30,
  30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30,
  28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158,
  28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158,
  28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158,
  28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158, 
    28.6842105263158, 28.6842105263158, 28.6842105263158, 28.6842105263158,
  27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316,
  27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316,
  27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316,
  27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316, 
    27.3684210526316, 27.3684210526316, 27.3684210526316, 27.3684210526316,
  26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474,
  26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474,
  26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474,
  26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474, 
    26.0526315789474, 26.0526315789474, 26.0526315789474, 26.0526315789474,
  24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632,
  24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632,
  24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632,
  24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632, 
    24.7368421052632, 24.7368421052632, 24.7368421052632, 24.7368421052632,
  23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789,
  23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789,
  23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789,
  23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789, 
    23.4210526315789, 23.4210526315789, 23.4210526315789, 23.4210526315789,
  22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947,
  22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947,
  22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947,
  22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947, 
    22.1052631578947, 22.1052631578947, 22.1052631578947, 22.1052631578947,
  20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105,
  20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105,
  20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105,
  20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105, 
    20.7894736842105, 20.7894736842105, 20.7894736842105, 20.7894736842105,
  19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263,
  19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263,
  19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263,
  19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263, 
    19.4736842105263, 19.4736842105263, 19.4736842105263, 19.4736842105263,
  18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421,
  18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421,
  18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421,
  18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421, 
    18.1578947368421, 18.1578947368421, 18.1578947368421, 18.1578947368421,
  16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579,
  16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579,
  16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579,
  16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579, 
    16.8421052631579, 16.8421052631579, 16.8421052631579, 16.8421052631579,
  15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737,
  15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737,
  15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737,
  15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737, 
    15.5263157894737, 15.5263157894737, 15.5263157894737, 15.5263157894737,
  14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895,
  14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895,
  14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895,
  14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895, 
    14.2105263157895, 14.2105263157895, 14.2105263157895, 14.2105263157895,
  12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053,
  12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053,
  12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053,
  12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053, 
    12.8947368421053, 12.8947368421053, 12.8947368421053, 12.8947368421053,
  11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211,
  11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211,
  11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211,
  11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211, 
    11.5789473684211, 11.5789473684211, 11.5789473684211, 11.5789473684211,
  10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368,
  10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368,
  10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368,
  10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368, 
    10.2631578947368, 10.2631578947368, 10.2631578947368, 10.2631578947368,
  8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263,
  8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263,
  8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263,
  8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263, 
    8.94736842105263, 8.94736842105263, 8.94736842105263, 8.94736842105263,
  7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842,
  7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842,
  7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842,
  7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842, 
    7.63157894736842, 7.63157894736842, 7.63157894736842, 7.63157894736842,
  6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421,
  6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421,
  6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421,
  6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421, 
    6.31578947368421, 6.31578947368421, 6.31578947368421, 6.31578947368421,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5 ;

 salt =
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35 ;

 h =
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001,
  19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001,
  19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001,
  19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001,
  19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 19.9981, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001 ;
}
