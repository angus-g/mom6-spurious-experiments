netcdf input_rho {
dimensions:
	x = 50 ;
	y = 4 ;
	z = 20 ;
variables:
	double x(x) ;
		x:_FillValue = NaN ;
	double y(y) ;
		y:_FillValue = NaN ;
	double z(z) ;
		z:_FillValue = NaN ;
	double temp(z, y, x) ;
		temp:_FillValue = NaN ;
	double salt(z, y, x) ;
		salt:_FillValue = NaN ;
	double h(z, y, x) ;
		h:_FillValue = NaN ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
data:

 x = 2.5, 7.5, 12.5, 17.5, 22.5, 27.5, 32.5, 37.5, 42.5, 47.5, 52.5, 57.5, 
    62.5, 67.5, 72.5, 77.5, 82.5, 87.5, 92.5, 97.5, 102.5, 107.5, 112.5, 
    117.5, 122.5, 127.5, 132.5, 137.5, 142.5, 147.5, 152.5, 157.5, 162.5, 
    167.5, 172.5, 177.5, 182.5, 187.5, 192.5, 197.5, 202.5, 207.5, 212.5, 
    217.5, 222.5, 227.5, 232.5, 237.5, 242.5, 247.5 ;

 y = 0, 1, 2, 3 ;

 z = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19 ;

 temp =
  19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75,
  19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75,
  19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75,
  19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 
    19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75, 19.75,
  19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25,
  19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25,
  19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25,
  19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 
    19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25, 19.25,
  18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75,
  18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75,
  18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75,
  18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 
    18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75, 18.75,
  18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25,
  18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25,
  18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25,
  18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 
    18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25, 18.25,
  17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75,
  17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75,
  17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75,
  17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 
    17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75, 17.75,
  17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25,
  17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25,
  17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25,
  17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 
    17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25, 17.25,
  16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75,
  16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75,
  16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75,
  16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 
    16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75, 16.75,
  16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25,
  16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25,
  16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25,
  16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 
    16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25, 16.25,
  15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75,
  15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75,
  15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75,
  15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 
    15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75, 15.75,
  15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25,
  15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25,
  15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25,
  15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 
    15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25, 15.25,
  14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75,
  14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75,
  14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75,
  14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 
    14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75, 14.75,
  14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25,
  14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25,
  14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25,
  14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 
    14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25, 14.25,
  13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75,
  13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75,
  13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75,
  13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 
    13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75, 13.75,
  13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25,
  13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25,
  13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25,
  13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 
    13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25, 13.25,
  12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75,
  12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75,
  12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75,
  12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 
    12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75, 12.75,
  12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25,
  12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25,
  12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25,
  12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 
    12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25, 12.25,
  11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75,
  11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75,
  11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75,
  11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 
    11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75, 11.75,
  11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25,
  11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25,
  11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25,
  11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 
    11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25, 11.25,
  10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75,
  10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75,
  10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75,
  10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 
    10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75, 10.75,
  10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25,
  10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25,
  10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25,
  10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 
    10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25, 10.25 ;

 salt =
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35 ;

 h =
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.8296469307822, 21.8108336932724, 20.1644723160189, 18.8319660892447, 
    17.7656073084617, 16.927612874677, 16.2888220020048, 15.8274499642497, 
    15.5280543733149, 15.380762217786, 15.380762217786, 15.5280543733149, 
    15.8274499642497, 16.2888220020048, 16.927612874677, 17.7656073084617, 
    18.8319660892447, 20.1644723160189, 21.8108336932724, 23.8296469307822, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.8296469307822, 21.8108336932724, 20.1644723160189, 18.8319660892447, 
    17.7656073084617, 16.927612874677, 16.2888220020048, 15.8274499642497, 
    15.5280543733149, 15.380762217786, 15.380762217786, 15.5280543733149, 
    15.8274499642497, 16.2888220020048, 16.927612874677, 17.7656073084617, 
    18.8319660892447, 20.1644723160189, 21.8108336932724, 23.8296469307822, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.8296469307822, 21.8108336932724, 20.1644723160189, 18.8319660892447, 
    17.7656073084617, 16.927612874677, 16.2888220020048, 15.8274499642497, 
    15.5280543733149, 15.380762217786, 15.380762217786, 15.5280543733149, 
    15.8274499642497, 16.2888220020048, 16.927612874677, 17.7656073084617, 
    18.8319660892447, 20.1644723160189, 21.8108336932724, 23.8296469307822, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.8296469307822, 21.8108336932724, 20.1644723160189, 18.8319660892447, 
    17.7656073084617, 16.927612874677, 16.2888220020048, 15.8274499642497, 
    15.5280543733149, 15.380762217786, 15.380762217786, 15.5280543733149, 
    15.8274499642497, 16.2888220020048, 16.927612874677, 17.7656073084617, 
    18.8319660892447, 20.1644723160189, 21.8108336932724, 23.8296469307822, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.8546567893742, 21.8632348876541, 20.2273532277594, 18.8973549140223, 
    17.8300227681635, 16.9898023605393, 16.3486221515312, 15.8852174768344, 
    15.5843853167429, 15.4363561048899, 15.4363561048899, 15.5843853167429, 
    15.8852174768344, 16.3486221515312, 16.9898023605393, 17.8300227681635, 
    18.8973549140223, 20.2273532277594, 21.8632348876541, 23.8546567893742, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.8546567893742, 21.8632348876541, 20.2273532277594, 18.8973549140223, 
    17.8300227681635, 16.9898023605393, 16.3486221515312, 15.8852174768344, 
    15.5843853167429, 15.4363561048899, 15.4363561048899, 15.5843853167429, 
    15.8852174768344, 16.3486221515312, 16.9898023605393, 17.8300227681635, 
    18.8973549140223, 20.2273532277594, 21.8632348876541, 23.8546567893742, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.8546567893742, 21.8632348876541, 20.2273532277594, 18.8973549140223, 
    17.8300227681635, 16.9898023605393, 16.3486221515312, 15.8852174768344, 
    15.5843853167429, 15.4363561048899, 15.4363561048899, 15.5843853167429, 
    15.8852174768344, 16.3486221515312, 16.9898023605393, 17.8300227681635, 
    18.8973549140223, 20.2273532277594, 21.8632348876541, 23.8546567893742, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.8546567893742, 21.8632348876541, 20.2273532277594, 18.8973549140223, 
    17.8300227681635, 16.9898023605393, 16.3486221515312, 15.8852174768344, 
    15.5843853167429, 15.4363561048899, 15.4363561048899, 15.5843853167429, 
    15.8852174768344, 16.3486221515312, 16.9898023605393, 17.8300227681635, 
    18.8973549140223, 20.2273532277594, 21.8632348876541, 23.8546567893742, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.904374236129, 21.9683014880961, 20.354061090677, 19.0294894571202, 
    17.9603940139917, 17.1157730021004, 16.469803413392, 16.0023021914225, 
    15.6985672857748, 15.5490469551031, 15.5490469551031, 15.6985672857748, 
    16.0023021914225, 16.469803413392, 17.1157730021004, 17.9603940139917, 
    19.0294894571202, 20.354061090677, 21.9683014880961, 23.904374236129, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.904374236129, 21.9683014880961, 20.354061090677, 19.0294894571202, 
    17.9603940139917, 17.1157730021004, 16.469803413392, 16.0023021914225, 
    15.6985672857748, 15.5490469551031, 15.5490469551031, 15.6985672857748, 
    16.0023021914225, 16.469803413392, 17.1157730021004, 17.9603940139917, 
    19.0294894571202, 20.354061090677, 21.9683014880961, 23.904374236129, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.904374236129, 21.9683014880961, 20.354061090677, 19.0294894571202, 
    17.9603940139917, 17.1157730021004, 16.469803413392, 16.0023021914225, 
    15.6985672857748, 15.5490469551031, 15.5490469551031, 15.6985672857748, 
    16.0023021914225, 16.469803413392, 17.1157730021004, 17.9603940139917, 
    19.0294894571202, 20.354061090677, 21.9683014880961, 23.904374236129, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.904374236129, 21.9683014880961, 20.354061090677, 19.0294894571202, 
    17.9603940139917, 17.1157730021004, 16.469803413392, 16.0023021914225, 
    15.6985672857748, 15.5490469551031, 15.5490469551031, 15.6985672857748, 
    16.0023021914225, 16.469803413392, 17.1157730021004, 17.9603940139917, 
    19.0294894571202, 20.354061090677, 21.9683014880961, 23.904374236129, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.9781822095507, 22.1265308814271, 20.5464970171389, 19.2311384432758, 
    18.1598868746678, 17.3088085284825, 16.6556339312114, 16.1819108934963, 
    15.8737473647065, 15.7219472628971, 15.7219472628971, 15.8737473647065, 
    16.1819108934963, 16.6556339312114, 17.3088085284825, 18.1598868746678, 
    19.2311384432758, 20.5464970171389, 22.1265308814271, 23.9781822095507, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.9781822095507, 22.1265308814271, 20.5464970171389, 19.2311384432758, 
    18.1598868746678, 17.3088085284825, 16.6556339312114, 16.1819108934963, 
    15.8737473647065, 15.7219472628971, 15.7219472628971, 15.8737473647065, 
    16.1819108934963, 16.6556339312114, 17.3088085284825, 18.1598868746678, 
    19.2311384432758, 20.5464970171389, 22.1265308814271, 23.9781822095507, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.9781822095507, 22.1265308814271, 20.5464970171389, 19.2311384432758, 
    18.1598868746678, 17.3088085284825, 16.6556339312114, 16.1819108934963, 
    15.8737473647065, 15.7219472628971, 15.7219472628971, 15.8737473647065, 
    16.1819108934963, 16.6556339312114, 17.3088085284825, 18.1598868746678, 
    19.2311384432758, 20.5464970171389, 22.1265308814271, 23.9781822095507, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    23.9781822095507, 22.1265308814271, 20.5464970171389, 19.2311384432758, 
    18.1598868746678, 17.3088085284825, 16.6556339312114, 16.1819108934963, 
    15.8737473647065, 15.7219472628971, 15.7219472628971, 15.8737473647065, 
    16.1819108934963, 16.6556339312114, 17.3088085284825, 18.1598868746678, 
    19.2311384432758, 20.5464970171389, 22.1265308814271, 23.9781822095507, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.0751244294751, 22.3385869245099, 20.8075307891426, 19.5065937604535, 
    18.4334703923934, 17.5740966936817, 16.9112946250701, 16.4291362735452, 
    16.1149277528913, 15.9600059617427, 15.9600059617427, 16.1149277528913, 
    16.4291362735452, 16.9112946250701, 17.5740966936817, 18.4334703923934, 
    19.5065937604535, 20.8075307891426, 22.3385869245099, 24.0751244294751, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.0751244294751, 22.3385869245099, 20.8075307891426, 19.5065937604535, 
    18.4334703923934, 17.5740966936817, 16.9112946250701, 16.4291362735452, 
    16.1149277528913, 15.9600059617427, 15.9600059617427, 16.1149277528913, 
    16.4291362735452, 16.9112946250701, 17.5740966936817, 18.4334703923934, 
    19.5065937604535, 20.8075307891426, 22.3385869245099, 24.0751244294751, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.0751244294751, 22.3385869245099, 20.8075307891426, 19.5065937604535, 
    18.4334703923934, 17.5740966936817, 16.9112946250701, 16.4291362735452, 
    16.1149277528913, 15.9600059617427, 15.9600059617427, 16.1149277528913, 
    16.4291362735452, 16.9112946250701, 17.5740966936817, 18.4334703923934, 
    19.5065937604535, 20.8075307891426, 22.3385869245099, 24.0751244294751, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.0751244294751, 22.3385869245099, 20.8075307891426, 19.5065937604535, 
    18.4334703923934, 17.5740966936817, 16.9112946250701, 16.4291362735452, 
    16.1149277528913, 15.9600059617427, 15.9600059617427, 16.1149277528913, 
    16.4291362735452, 16.9112946250701, 17.5740966936817, 18.4334703923934, 
    19.5065937604535, 20.8075307891426, 22.3385869245099, 24.0751244294751, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.1938704098673, 22.6051879930684, 21.1410086316465, 19.8618402636631, 
    18.7882023737792, 17.9190769868436, 17.2442530246281, 16.7513380516875, 
    16.429346706479, 16.2703879425722, 16.2703879425722, 16.429346706479, 
    16.7513380516875, 17.2442530246281, 17.9190769868436, 18.7882023737792, 
    19.8618402636631, 21.1410086316465, 22.6051879930684, 24.1938704098673, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.1938704098673, 22.6051879930684, 21.1410086316465, 19.8618402636631, 
    18.7882023737792, 17.9190769868436, 17.2442530246281, 16.7513380516875, 
    16.429346706479, 16.2703879425722, 16.2703879425722, 16.429346706479, 
    16.7513380516875, 17.2442530246281, 17.9190769868436, 18.7882023737792, 
    19.8618402636631, 21.1410086316465, 22.6051879930684, 24.1938704098673, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.1938704098673, 22.6051879930684, 21.1410086316465, 19.8618402636631, 
    18.7882023737792, 17.9190769868436, 17.2442530246281, 16.7513380516875, 
    16.429346706479, 16.2703879425722, 16.2703879425722, 16.429346706479, 
    16.7513380516875, 17.2442530246281, 17.9190769868436, 18.7882023737792, 
    19.8618402636631, 21.1410086316465, 22.6051879930684, 24.1938704098673, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.1938704098673, 22.6051879930684, 21.1410086316465, 19.8618402636631, 
    18.7882023737792, 17.9190769868436, 17.2442530246281, 16.7513380516875, 
    16.429346706479, 16.2703879425722, 16.2703879425722, 16.429346706479, 
    16.7513380516875, 17.2442530246281, 17.9190769868436, 18.7882023737792, 
    19.8618402636631, 21.1410086316465, 22.6051879930684, 24.1938704098673, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.3326722241113, 22.9269347466473, 21.5517356025668, 20.3047845454261, 
    19.2336470410445, 18.3539651485402, 17.6648356572618, 17.1587309761422, 
    16.82706847192, 16.6630626966011, 16.6630626966011, 16.82706847192, 
    17.1587309761422, 17.6648356572618, 18.3539651485402, 19.2336470410445, 
    20.3047845454261, 21.5517356025668, 22.9269347466473, 24.3326722241113, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.3326722241113, 22.9269347466473, 21.5517356025668, 20.3047845454261, 
    19.2336470410445, 18.3539651485402, 17.6648356572618, 17.1587309761422, 
    16.82706847192, 16.6630626966011, 16.6630626966011, 16.82706847192, 
    17.1587309761422, 17.6648356572618, 18.3539651485402, 19.2336470410445, 
    20.3047845454261, 21.5517356025668, 22.9269347466473, 24.3326722241113, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.3326722241113, 22.9269347466473, 21.5517356025668, 20.3047845454261, 
    19.2336470410445, 18.3539651485402, 17.6648356572618, 17.1587309761422, 
    16.82706847192, 16.6630626966011, 16.6630626966011, 16.82706847192, 
    17.1587309761422, 17.6648356572618, 18.3539651485402, 19.2336470410445, 
    20.3047845454261, 21.5517356025668, 22.9269347466473, 24.3326722241113, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.3326722241113, 22.9269347466473, 21.5517356025668, 20.3047845454261, 
    19.2336470410445, 18.3539651485402, 17.6648356572618, 17.1587309761422, 
    16.82706847192, 16.6630626966011, 16.6630626966011, 16.82706847192, 
    17.1587309761422, 17.6648356572618, 18.3539651485402, 19.2336470410445, 
    20.3047845454261, 21.5517356025668, 22.9269347466473, 24.3326722241113, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.4893166189955, 23.304056687434, 22.0453980243628, 20.8455366725627, 
    19.7824588918212, 18.8925191167478, 18.1870813083334, 17.6652705519531, 
    17.3218765418669, 17.1516975244433, 17.1516975244433, 17.3218765418669, 
    17.6652705519531, 18.1870813083334, 18.8925191167478, 19.7824588918212, 
    20.8455366725627, 22.0453980243628, 23.304056687434, 24.4893166189955, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.4893166189955, 23.304056687434, 22.0453980243628, 20.8455366725627, 
    19.7824588918212, 18.8925191167478, 18.1870813083334, 17.6652705519531, 
    17.3218765418669, 17.1516975244433, 17.1516975244433, 17.3218765418669, 
    17.6652705519531, 18.1870813083334, 18.8925191167478, 19.7824588918212, 
    20.8455366725627, 22.0453980243628, 23.304056687434, 24.4893166189955, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.4893166189955, 23.304056687434, 22.0453980243628, 20.8455366725627, 
    19.7824588918212, 18.8925191167478, 18.1870813083334, 17.6652705519531, 
    17.3218765418669, 17.1516975244433, 17.1516975244433, 17.3218765418669, 
    17.6652705519531, 18.1870813083334, 18.8925191167478, 19.7824588918212, 
    20.8455366725627, 22.0453980243628, 23.304056687434, 24.4893166189955, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.4893166189955, 23.304056687434, 22.0453980243628, 20.8455366725627, 
    19.7824588918212, 18.8925191167478, 18.1870813083334, 17.6652705519531, 
    17.3218765418669, 17.1516975244433, 17.1516975244433, 17.3218765418669, 
    17.6652705519531, 18.1870813083334, 18.8925191167478, 19.7824588918212, 
    20.8455366725627, 22.0453980243628, 23.304056687434, 24.4893166189955, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.6610777172359, 23.7360509964541, 22.6283667279538, 21.4967219198757, 
    20.4511759038873, 19.5531448833227, 18.8300077404276, 18.2899864804067, 
    17.9326277737055, 17.7550154668227, 17.7550154668227, 17.9326277737055, 
    18.2899864804067, 18.8300077404276, 19.5531448833227, 20.4511759038873, 
    21.4967219198757, 22.6283667279538, 23.7360509964541, 24.6610777172359, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.6610777172359, 23.7360509964541, 22.6283667279538, 21.4967219198757, 
    20.4511759038873, 19.5531448833227, 18.8300077404276, 18.2899864804067, 
    17.9326277737055, 17.7550154668227, 17.7550154668227, 17.9326277737055, 
    18.2899864804067, 18.8300077404276, 19.5531448833227, 20.4511759038873, 
    21.4967219198757, 22.6283667279538, 23.7360509964541, 24.6610777172359, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.6610777172359, 23.7360509964541, 22.6283667279538, 21.4967219198757, 
    20.4511759038873, 19.5531448833227, 18.8300077404276, 18.2899864804067, 
    17.9326277737055, 17.7550154668227, 17.7550154668227, 17.9326277737055, 
    18.2899864804067, 18.8300077404276, 19.5531448833227, 20.4511759038873, 
    21.4967219198757, 22.6283667279538, 23.7360509964541, 24.6610777172359, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.6610777172359, 23.7360509964541, 22.6283667279538, 21.4967219198757, 
    20.4511759038873, 19.5531448833227, 18.8300077404276, 18.2899864804067, 
    17.9326277737055, 17.7550154668227, 17.7550154668227, 17.9326277737055, 
    18.2899864804067, 18.8300077404276, 19.5531448833227, 20.4511759038873, 
    21.4967219198757, 22.6283667279538, 23.7360509964541, 24.6610777172359, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.8446775058025, 24.2211837404477, 23.3072822931047, 22.273760738328, 
    21.2612673517159, 20.3604890316332, 19.6195058682658, 19.0590141307703, 
    18.685334450637, 18.4988911958477, 18.4988911958477, 18.685334450637, 
    19.0590141307703, 19.6195058682658, 20.3604890316332, 21.2612673517159, 
    22.273760738328, 23.3072822931047, 24.2211837404477, 24.8446775058025, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.8446775058025, 24.2211837404477, 23.3072822931047, 22.273760738328, 
    21.2612673517159, 20.3604890316332, 19.6195058682658, 19.0590141307703, 
    18.685334450637, 18.4988911958477, 18.4988911958477, 18.685334450637, 
    19.0590141307703, 19.6195058682658, 20.3604890316332, 21.2612673517159, 
    22.273760738328, 23.3072822931047, 24.2211837404477, 24.8446775058025, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.8446775058025, 24.2211837404477, 23.3072822931047, 22.273760738328, 
    21.2612673517159, 20.3604890316332, 19.6195058682658, 19.0590141307703, 
    18.685334450637, 18.4988911958477, 18.4988911958477, 18.685334450637, 
    19.0590141307703, 19.6195058682658, 20.3604890316332, 21.2612673517159, 
    22.273760738328, 23.3072822931047, 24.2211837404477, 24.8446775058025, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    24.8446775058025, 24.2211837404477, 23.3072822931047, 22.273760738328, 
    21.2612673517159, 20.3604890316332, 19.6195058682658, 19.0590141307703, 
    18.685334450637, 18.4988911958477, 18.4988911958477, 18.685334450637, 
    19.0590141307703, 19.6195058682658, 20.3604890316332, 21.2612673517159, 
    22.273760738328, 23.3072822931047, 24.2211837404477, 24.8446775058025, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25.03626339557, 
    24.7558263516493, 24.0882627313388, 23.1949718399376, 22.2404590991992, 
    21.3477294185654, 20.5912091449121, 20.0087501797549, 19.6164386499739, 
    19.4196639890118, 19.4196639890118, 19.6164386499739, 20.0087501797549, 
    20.5912091449121, 21.3477294185654, 22.2404590991992, 23.1949718399376, 
    24.0882627313388, 24.7558263516493, 25.03626339557, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25.03626339557, 
    24.7558263516493, 24.0882627313388, 23.1949718399376, 22.2404590991992, 
    21.3477294185654, 20.5912091449121, 20.0087501797549, 19.6164386499739, 
    19.4196639890118, 19.4196639890118, 19.6164386499739, 20.0087501797549, 
    20.5912091449121, 21.3477294185654, 22.2404590991992, 23.1949718399376, 
    24.0882627313388, 24.7558263516493, 25.03626339557, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25.03626339557, 
    24.7558263516493, 24.0882627313388, 23.1949718399376, 22.2404590991992, 
    21.3477294185654, 20.5912091449121, 20.0087501797549, 19.6164386499739, 
    19.4196639890118, 19.4196639890118, 19.6164386499739, 20.0087501797549, 
    20.5912091449121, 21.3477294185654, 22.2404590991992, 23.1949718399376, 
    24.0882627313388, 24.7558263516493, 25.03626339557, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25.03626339557, 
    24.7558263516493, 24.0882627313388, 23.1949718399376, 22.2404590991992, 
    21.3477294185654, 20.5912091449121, 20.0087501797549, 19.6164386499739, 
    19.4196639890118, 19.4196639890118, 19.6164386499739, 20.0087501797549, 
    20.5912091449121, 21.3477294185654, 22.2404590991992, 23.1949718399376, 
    24.0882627313388, 24.7558263516493, 25.03626339557, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.2314139839538, 25.3336164346724, 24.9754883933963, 24.2811813587252, 
    23.4242646943941, 22.559845375413, 21.7949043935673, 21.190874452582, 
    20.7781115500938, 20.5695369135359, 20.5695369135359, 20.7781115500938, 
    21.190874452582, 21.7949043935673, 22.559845375413, 23.4242646943941, 
    24.2811813587252, 24.9754883933963, 25.3336164346724, 25.2314139839538, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.2314139839538, 25.3336164346724, 24.9754883933963, 24.2811813587252, 
    23.4242646943941, 22.559845375413, 21.7949043935673, 21.190874452582, 
    20.7781115500938, 20.5695369135359, 20.5695369135359, 20.7781115500938, 
    21.190874452582, 21.7949043935673, 22.559845375413, 23.4242646943941, 
    24.2811813587252, 24.9754883933963, 25.3336164346724, 25.2314139839538, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.2314139839538, 25.3336164346724, 24.9754883933963, 24.2811813587252, 
    23.4242646943941, 22.559845375413, 21.7949043935673, 21.190874452582, 
    20.7781115500938, 20.5695369135359, 20.5695369135359, 20.7781115500938, 
    21.190874452582, 21.7949043935673, 22.559845375413, 23.4242646943941, 
    24.2811813587252, 24.9754883933963, 25.3336164346724, 25.2314139839538, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.2314139839538, 25.3336164346724, 24.9754883933963, 24.2811813587252, 
    23.4242646943941, 22.559845375413, 21.7949043935673, 21.190874452582, 
    20.7781115500938, 20.5695369135359, 20.5695369135359, 20.7781115500938, 
    21.190874452582, 21.7949043935673, 22.559845375413, 23.4242646943941, 
    24.2811813587252, 24.9754883933963, 25.3336164346724, 25.2314139839538, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.4251851613234, 25.944472338988, 25.9688177571947, 25.5541811742133, 
    24.857360063427, 24.0581602805123, 23.3013899627234, 22.6805557954933, 
    22.2471206521761, 22.0256996234475, 22.0256996234475, 22.2471206521761, 
    22.6805557954933, 23.3013899627234, 24.0581602805123, 24.857360063427, 
    25.5541811742133, 25.9688177571947, 25.944472338988, 25.4251851613234, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.4251851613234, 25.944472338988, 25.9688177571947, 25.5541811742133, 
    24.857360063427, 24.0581602805123, 23.3013899627234, 22.6805557954933, 
    22.2471206521761, 22.0256996234475, 22.0256996234475, 22.2471206521761, 
    22.6805557954933, 23.3013899627234, 24.0581602805123, 24.857360063427, 
    25.5541811742133, 25.9688177571947, 25.944472338988, 25.4251851613234, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.4251851613234, 25.944472338988, 25.9688177571947, 25.5541811742133, 
    24.857360063427, 24.0581602805123, 23.3013899627234, 22.6805557954933, 
    22.2471206521761, 22.0256996234475, 22.0256996234475, 22.2471206521761, 
    22.6805557954933, 23.3013899627234, 24.0581602805123, 24.857360063427, 
    25.5541811742133, 25.9688177571947, 25.944472338988, 25.4251851613234, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.4251851613234, 25.944472338988, 25.9688177571947, 25.5541811742133, 
    24.857360063427, 24.0581602805123, 23.3013899627234, 22.6805557954933, 
    22.2471206521761, 22.0256996234475, 22.0256996234475, 22.2471206521761, 
    22.6805557954933, 23.3013899627234, 24.0581602805123, 24.857360063427, 
    25.5541811742133, 25.9688177571947, 25.944472338988, 25.4251851613234, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.6122080865181, 26.5735685175113, 27.0600209209555, 27.0327502988659, 
    26.5936416166563, 25.9261519532193, 25.2131239428117, 24.5901961933143, 
    24.1402111642773, 23.9063799992776, 23.9063799992776, 24.1402111642773, 
    24.5901961933143, 25.2131239428117, 25.9261519532193, 26.5936416166563, 
    27.0327502988659, 27.0600209209555, 26.5735685175113, 25.6122080865181, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.6122080865181, 26.5735685175113, 27.0600209209555, 27.0327502988659, 
    26.5936416166563, 25.9261519532193, 25.2131239428117, 24.5901961933143, 
    24.1402111642773, 23.9063799992776, 23.9063799992776, 24.1402111642773, 
    24.5901961933143, 25.2131239428117, 25.9261519532193, 26.5936416166563, 
    27.0327502988659, 27.0600209209555, 26.5735685175113, 25.6122080865181, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.6122080865181, 26.5735685175113, 27.0600209209555, 27.0327502988659, 
    26.5936416166563, 25.9261519532193, 25.2131239428117, 24.5901961933143, 
    24.1402111642773, 23.9063799992776, 23.9063799992776, 24.1402111642773, 
    24.5901961933143, 25.2131239428117, 25.9261519532193, 26.5936416166563, 
    27.0327502988659, 27.0600209209555, 26.5735685175113, 25.6122080865181, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.6122080865181, 26.5735685175113, 27.0600209209555, 27.0327502988659, 
    26.5936416166563, 25.9261519532193, 25.2131239428117, 24.5901961933143, 
    24.1402111642773, 23.9063799992776, 23.9063799992776, 24.1402111642773, 
    24.5901961933143, 25.2131239428117, 25.9261519532193, 26.5936416166563, 
    27.0327502988659, 27.0600209209555, 26.5735685175113, 25.6122080865181, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.7868474736291, 27.2005011592135, 28.2273286839547, 28.7239322426845, 
    28.6917660667959, 28.2750357624696, 27.6801143330499, 27.092758625336, 
    26.6417056388756, 26.4002910793875, 26.4002910793875, 26.6417056388756, 
    27.092758625336, 27.6801143330499, 28.2750357624696, 28.6917660667959, 
    28.7239322426845, 28.2273286839547, 27.2005011592135, 25.7868474736291, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.7868474736291, 27.2005011592135, 28.2273286839547, 28.7239322426845, 
    28.6917660667959, 28.2750357624696, 27.6801143330499, 27.092758625336, 
    26.6417056388756, 26.4002910793875, 26.4002910793875, 26.6417056388756, 
    27.092758625336, 27.6801143330499, 28.2750357624696, 28.6917660667959, 
    28.7239322426845, 28.2273286839547, 27.2005011592135, 25.7868474736291, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.7868474736291, 27.2005011592135, 28.2273286839547, 28.7239322426845, 
    28.6917660667959, 28.2750357624696, 27.6801143330499, 27.092758625336, 
    26.6417056388756, 26.4002910793875, 26.4002910793875, 26.6417056388756, 
    27.092758625336, 27.6801143330499, 28.2750357624696, 28.6917660667959, 
    28.7239322426845, 28.2273286839547, 27.2005011592135, 25.7868474736291, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.7868474736291, 27.2005011592135, 28.2273286839547, 28.7239322426845, 
    28.6917660667959, 28.2750357624696, 27.6801143330499, 27.092758625336, 
    26.6417056388756, 26.4002910793875, 26.4002910793875, 26.6417056388756, 
    27.092758625336, 27.6801143330499, 28.2750357624696, 28.6917660667959, 
    28.7239322426845, 28.2273286839547, 27.2005011592135, 25.7868474736291, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.9434224613103, 27.7990263700528, 29.4285894216251, 30.6061005930228, 
    31.1982021080483, 31.2420125761087, 30.9198569249714, 30.4602765469147, 
    30.0538627187645, 29.8224422621923, 29.8224422621923, 30.0538627187645, 
    30.4602765469147, 30.9198569249714, 31.2420125761087, 31.1982021080483, 
    30.6061005930228, 29.4285894216251, 27.7990263700528, 25.9434224613103, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.9434224613103, 27.7990263700528, 29.4285894216251, 30.6061005930228, 
    31.1982021080483, 31.2420125761087, 30.9198569249714, 30.4602765469147, 
    30.0538627187645, 29.8224422621923, 29.8224422621923, 30.0538627187645, 
    30.4602765469147, 30.9198569249714, 31.2420125761087, 31.1982021080483, 
    30.6061005930228, 29.4285894216251, 27.7990263700528, 25.9434224613103, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.9434224613103, 27.7990263700528, 29.4285894216251, 30.6061005930228, 
    31.1982021080483, 31.2420125761087, 30.9198569249714, 30.4602765469147, 
    30.0538627187645, 29.8224422621923, 29.8224422621923, 30.0538627187645, 
    30.4602765469147, 30.9198569249714, 31.2420125761087, 31.1982021080483, 
    30.6061005930228, 29.4285894216251, 27.7990263700528, 25.9434224613103, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25.9434224613103, 27.7990263700528, 29.4285894216251, 30.6061005930228, 
    31.1982021080483, 31.2420125761087, 30.9198569249714, 30.4602765469147, 
    30.0538627187645, 29.8224422621923, 29.8224422621923, 30.0538627187645, 
    30.4602765469147, 30.9198569249714, 31.2420125761087, 31.1982021080483, 
    30.6061005930228, 29.4285894216251, 27.7990263700528, 25.9434224613103, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.0764830767929, 28.3378742052888, 30.5948411856911, 32.600741534627, 
    34.1007231334441, 34.9556579816398, 35.2232161157257, 35.1160327966077, 
    34.883640170719, 34.7182333298409, 34.7182333298409, 34.883640170719, 
    35.1160327966077, 35.2232161157257, 34.9556579816398, 34.1007231334441, 
    32.600741534627, 30.5948411856911, 28.3378742052888, 26.0764830767929, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.0764830767929, 28.3378742052888, 30.5948411856911, 32.600741534627, 
    34.1007231334441, 34.9556579816398, 35.2232161157257, 35.1160327966077, 
    34.883640170719, 34.7182333298409, 34.7182333298409, 34.883640170719, 
    35.1160327966077, 35.2232161157257, 34.9556579816398, 34.1007231334441, 
    32.600741534627, 30.5948411856911, 28.3378742052888, 26.0764830767929, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.0764830767929, 28.3378742052888, 30.5948411856911, 32.600741534627, 
    34.1007231334441, 34.9556579816398, 35.2232161157257, 35.1160327966077, 
    34.883640170719, 34.7182333298409, 34.7182333298409, 34.883640170719, 
    35.1160327966077, 35.2232161157257, 34.9556579816398, 34.1007231334441, 
    32.600741534627, 30.5948411856911, 28.3378742052888, 26.0764830767929, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.0764830767929, 28.3378742052888, 30.5948411856911, 32.600741534627, 
    34.1007231334441, 34.9556579816398, 35.2232161157257, 35.1160327966077, 
    34.883640170719, 34.7182333298409, 34.7182333298409, 34.883640170719, 
    35.1160327966077, 35.2232161157257, 34.9556579816398, 34.1007231334441, 
    32.600741534627, 30.5948411856911, 28.3378742052888, 26.0764830767929, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.1811239729895, 28.7831067799539, 31.6286591500135, 34.5370015581166, 
    37.2273246489354, 39.3941639251915, 40.8500207562171, 41.626399836289, 
    41.9317080024242, 42.0088607293264, 42.0088607293264, 41.9317080024242, 
    41.626399836289, 40.8500207562171, 39.3941639251915, 37.2273246489354, 
    34.5370015581166, 31.6286591500135, 28.7831067799539, 26.1811239729895, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.1811239729895, 28.7831067799539, 31.6286591500135, 34.5370015581166, 
    37.2273246489354, 39.3941639251915, 40.8500207562171, 41.626399836289, 
    41.9317080024242, 42.0088607293264, 42.0088607293264, 41.9317080024242, 
    41.626399836289, 40.8500207562171, 39.3941639251915, 37.2273246489354, 
    34.5370015581166, 31.6286591500135, 28.7831067799539, 26.1811239729895, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.1811239729895, 28.7831067799539, 31.6286591500135, 34.5370015581166, 
    37.2273246489354, 39.3941639251915, 40.8500207562171, 41.626399836289, 
    41.9317080024242, 42.0088607293264, 42.0088607293264, 41.9317080024242, 
    41.626399836289, 40.8500207562171, 39.3941639251915, 37.2273246489354, 
    34.5370015581166, 31.6286591500135, 28.7831067799539, 26.1811239729895, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.1811239729895, 28.7831067799539, 31.6286591500135, 34.5370015581166, 
    37.2273246489354, 39.3941639251915, 40.8500207562171, 41.626399836289, 
    41.9317080024242, 42.0088607293264, 42.0088607293264, 41.9317080024242, 
    41.626399836289, 40.8500207562171, 39.3941639251915, 37.2273246489354, 
    34.5370015581166, 31.6286591500135, 28.7831067799539, 26.1811239729895, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.2533059059365, 29.1021505760053, 32.4138028255732, 36.1343879579156, 
    40.0986339154295, 44.0055096597119, 47.4660784282842, 50.1408072898158, 
    51.8755709333527, 52.7022506428348, 52.7022506428348, 51.8755709333527, 
    50.1408072898158, 47.4660784282842, 44.0055096597119, 40.0986339154295, 
    36.1343879579156, 32.4138028255732, 29.1021505760053, 26.2533059059365, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.2533059059365, 29.1021505760053, 32.4138028255732, 36.1343879579156, 
    40.0986339154295, 44.0055096597119, 47.4660784282842, 50.1408072898158, 
    51.8755709333527, 52.7022506428348, 52.7022506428348, 51.8755709333527, 
    50.1408072898158, 47.4660784282842, 44.0055096597119, 40.0986339154295, 
    36.1343879579156, 32.4138028255732, 29.1021505760053, 26.2533059059365, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.2533059059365, 29.1021505760053, 32.4138028255732, 36.1343879579156, 
    40.0986339154295, 44.0055096597119, 47.4660784282842, 50.1408072898158, 
    51.8755709333527, 52.7022506428348, 52.7022506428348, 51.8755709333527, 
    50.1408072898158, 47.4660784282842, 44.0055096597119, 40.0986339154295, 
    36.1343879579156, 32.4138028255732, 29.1021505760053, 26.2533059059365, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.2533059059365, 29.1021505760053, 32.4138028255732, 36.1343879579156, 
    40.0986339154295, 44.0055096597119, 47.4660784282842, 50.1408072898158, 
    51.8755709333527, 52.7022506428348, 52.7022506428348, 51.8755709333527, 
    50.1408072898158, 47.4660784282842, 44.0055096597119, 40.0986339154295, 
    36.1343879579156, 32.4138028255732, 29.1021505760053, 26.2533059059365, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.2901474106526, 29.2689552276536, 32.8404832098856, 37.0555646379193, 
    41.901491733744, 47.2404444406001, 52.740226275611, 57.8429912933845, 
    61.835694481304, 64.0394681024395, 64.0394681024395, 61.835694481304, 
    57.8429912933845, 52.740226275611, 47.2404444406001, 41.901491733744, 
    37.0555646379193, 32.8404832098856, 29.2689552276536, 26.2901474106526, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.2901474106526, 29.2689552276536, 32.8404832098856, 37.0555646379193, 
    41.901491733744, 47.2404444406001, 52.740226275611, 57.8429912933845, 
    61.835694481304, 64.0394681024395, 64.0394681024395, 61.835694481304, 
    57.8429912933845, 52.740226275611, 47.2404444406001, 41.901491733744, 
    37.0555646379193, 32.8404832098856, 29.2689552276536, 26.2901474106526, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.2901474106526, 29.2689552276536, 32.8404832098856, 37.0555646379193, 
    41.901491733744, 47.2404444406001, 52.740226275611, 57.8429912933845, 
    61.835694481304, 64.0394681024395, 64.0394681024395, 61.835694481304, 
    57.8429912933845, 52.740226275611, 47.2404444406001, 41.901491733744, 
    37.0555646379193, 32.8404832098856, 29.2689552276536, 26.2901474106526, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25,
  25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    26.2901474106526, 29.2689552276536, 32.8404832098856, 37.0555646379193, 
    41.901491733744, 47.2404444406001, 52.740226275611, 57.8429912933845, 
    61.835694481304, 64.0394681024395, 64.0394681024395, 61.835694481304, 
    57.8429912933845, 52.740226275611, 47.2404444406001, 41.901491733744, 
    37.0555646379193, 32.8404832098856, 29.2689552276536, 26.2901474106526, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25 ;
}
