netcdf input {
dimensions:
	x = 50 ;
	y = 4 ;
	z = 20 ;
variables:
	double x(x) ;
		x:_FillValue = NaN ;
	double y(y) ;
		y:_FillValue = NaN ;
	double z(z) ;
		z:_FillValue = NaN ;
	double temp(z, y, x) ;
		temp:_FillValue = NaN ;
	double salt(z, y, x) ;
		salt:_FillValue = NaN ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
data:

 x = 2.5, 7.5, 12.5, 17.5, 22.5, 27.5, 32.5, 37.5, 42.5, 47.5, 52.5, 57.5, 
    62.5, 67.5, 72.5, 77.5, 82.5, 87.5, 92.5, 97.5, 102.5, 107.5, 112.5, 
    117.5, 122.5, 127.5, 132.5, 137.5, 142.5, 147.5, 152.5, 157.5, 162.5, 
    167.5, 172.5, 177.5, 182.5, 187.5, 192.5, 197.5, 202.5, 207.5, 212.5, 
    217.5, 222.5, 227.5, 232.5, 237.5, 242.5, 247.5 ;

 y = 2.5, 7.5, 12.5, 17.5 ;

 z = 12.5, 37.5, 62.5, 87.5, 112.5, 137.5, 162.5, 187.5, 212.5, 237.5, 262.5, 
    287.5, 312.5, 337.5, 362.5, 387.5, 412.5, 437.5, 462.5, 487.5 ;

 temp =
  19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 17.8435986117215, 
    17.8435968430093, 17.8435952708202, 17.8435938951544, 17.8435927160121, 
    17.8435917333933, 17.8435909472981, 17.8435903577267, 17.8435899646791, 
    17.8435897681552, 17.8435897681552, 17.8435899646791, 17.8435903577267, 
    17.8435909472981, 17.8435917333933, 17.8435927160121, 17.8435938951544, 
    17.8435952708202, 17.8435968430093, 17.8435986117215, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897,
  19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 17.8435986117215, 
    17.8435968430093, 17.8435952708202, 17.8435938951544, 17.8435927160121, 
    17.8435917333933, 17.8435909472981, 17.8435903577267, 17.8435899646791, 
    17.8435897681552, 17.8435897681552, 17.8435899646791, 17.8435903577267, 
    17.8435909472981, 17.8435917333933, 17.8435927160121, 17.8435938951544, 
    17.8435952708202, 17.8435968430093, 17.8435986117215, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897,
  19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 17.8435986117215, 
    17.8435968430093, 17.8435952708202, 17.8435938951544, 17.8435927160121, 
    17.8435917333933, 17.8435909472981, 17.8435903577267, 17.8435899646791, 
    17.8435897681552, 17.8435897681552, 17.8435899646791, 17.8435903577267, 
    17.8435909472981, 17.8435917333933, 17.8435927160121, 17.8435938951544, 
    17.8435952708202, 17.8435968430093, 17.8435986117215, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897,
  19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 17.8435986117215, 
    17.8435968430093, 17.8435952708202, 17.8435938951544, 17.8435927160121, 
    17.8435917333933, 17.8435909472981, 17.8435903577267, 17.8435899646791, 
    17.8435897681552, 17.8435897681552, 17.8435899646791, 17.8435903577267, 
    17.8435909472981, 17.8435917333933, 17.8435927160121, 17.8435938951544, 
    17.8435952708202, 17.8435968430093, 17.8435986117215, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897, 19.8435897435897, 19.8435897435897, 
    19.8435897435897, 19.8435897435897,
  19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 17.330778098901, 
    17.3307763301888, 17.3307747579997, 17.3307733823339, 17.3307722031916, 
    17.3307712205728, 17.3307704344776, 17.3307698449062, 17.3307694518586, 
    17.3307692553347, 17.3307692553347, 17.3307694518586, 17.3307698449062, 
    17.3307704344776, 17.3307712205728, 17.3307722031916, 17.3307733823339, 
    17.3307747579997, 17.3307763301888, 17.330778098901, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692,
  19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 17.330778098901, 
    17.3307763301888, 17.3307747579997, 17.3307733823339, 17.3307722031916, 
    17.3307712205728, 17.3307704344776, 17.3307698449062, 17.3307694518586, 
    17.3307692553347, 17.3307692553347, 17.3307694518586, 17.3307698449062, 
    17.3307704344776, 17.3307712205728, 17.3307722031916, 17.3307733823339, 
    17.3307747579997, 17.3307763301888, 17.330778098901, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692,
  19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 17.330778098901, 
    17.3307763301888, 17.3307747579997, 17.3307733823339, 17.3307722031916, 
    17.3307712205728, 17.3307704344776, 17.3307698449062, 17.3307694518586, 
    17.3307692553347, 17.3307692553347, 17.3307694518586, 17.3307698449062, 
    17.3307704344776, 17.3307712205728, 17.3307722031916, 17.3307733823339, 
    17.3307747579997, 17.3307763301888, 17.330778098901, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692,
  19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 17.330778098901, 
    17.3307763301888, 17.3307747579997, 17.3307733823339, 17.3307722031916, 
    17.3307712205728, 17.3307704344776, 17.3307698449062, 17.3307694518586, 
    17.3307692553347, 17.3307692553347, 17.3307694518586, 17.3307698449062, 
    17.3307704344776, 17.3307712205728, 17.3307722031916, 17.3307733823339, 
    17.3307747579997, 17.3307763301888, 17.330778098901, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692, 19.3307692307692, 19.3307692307692, 
    19.3307692307692, 19.3307692307692,
  18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 16.8179575860805, 
    16.8179558173683, 16.8179542451792, 16.8179528695134, 16.8179516903711, 
    16.8179507077523, 16.8179499216571, 16.8179493320857, 16.817948939038, 
    16.8179487425142, 16.8179487425142, 16.817948939038, 16.8179493320857, 
    16.8179499216571, 16.8179507077523, 16.8179516903711, 16.8179528695134, 
    16.8179542451792, 16.8179558173683, 16.8179575860805, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487,
  18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 16.8179575860805, 
    16.8179558173683, 16.8179542451792, 16.8179528695134, 16.8179516903711, 
    16.8179507077523, 16.8179499216571, 16.8179493320857, 16.817948939038, 
    16.8179487425142, 16.8179487425142, 16.817948939038, 16.8179493320857, 
    16.8179499216571, 16.8179507077523, 16.8179516903711, 16.8179528695134, 
    16.8179542451792, 16.8179558173683, 16.8179575860805, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487,
  18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 16.8179575860805, 
    16.8179558173683, 16.8179542451792, 16.8179528695134, 16.8179516903711, 
    16.8179507077523, 16.8179499216571, 16.8179493320857, 16.817948939038, 
    16.8179487425142, 16.8179487425142, 16.817948939038, 16.8179493320857, 
    16.8179499216571, 16.8179507077523, 16.8179516903711, 16.8179528695134, 
    16.8179542451792, 16.8179558173683, 16.8179575860805, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487,
  18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 16.8179575860805, 
    16.8179558173683, 16.8179542451792, 16.8179528695134, 16.8179516903711, 
    16.8179507077523, 16.8179499216571, 16.8179493320857, 16.817948939038, 
    16.8179487425142, 16.8179487425142, 16.817948939038, 16.8179493320857, 
    16.8179499216571, 16.8179507077523, 16.8179516903711, 16.8179528695134, 
    16.8179542451792, 16.8179558173683, 16.8179575860805, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487, 18.8179487179487, 18.8179487179487, 
    18.8179487179487, 18.8179487179487,
  18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 16.3051370732599, 
    16.3051353045477, 16.3051337323587, 16.3051323566929, 16.3051311775506, 
    16.3051301949318, 16.3051294088366, 16.3051288192652, 16.3051284262175, 
    16.3051282296937, 16.3051282296937, 16.3051284262175, 16.3051288192652, 
    16.3051294088366, 16.3051301949318, 16.3051311775506, 16.3051323566929, 
    16.3051337323587, 16.3051353045477, 16.3051370732599, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282,
  18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 16.3051370732599, 
    16.3051353045477, 16.3051337323587, 16.3051323566929, 16.3051311775506, 
    16.3051301949318, 16.3051294088366, 16.3051288192652, 16.3051284262175, 
    16.3051282296937, 16.3051282296937, 16.3051284262175, 16.3051288192652, 
    16.3051294088366, 16.3051301949318, 16.3051311775506, 16.3051323566929, 
    16.3051337323587, 16.3051353045477, 16.3051370732599, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282,
  18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 16.3051370732599, 
    16.3051353045477, 16.3051337323587, 16.3051323566929, 16.3051311775506, 
    16.3051301949318, 16.3051294088366, 16.3051288192652, 16.3051284262175, 
    16.3051282296937, 16.3051282296937, 16.3051284262175, 16.3051288192652, 
    16.3051294088366, 16.3051301949318, 16.3051311775506, 16.3051323566929, 
    16.3051337323587, 16.3051353045477, 16.3051370732599, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282,
  18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 16.3051370732599, 
    16.3051353045477, 16.3051337323587, 16.3051323566929, 16.3051311775506, 
    16.3051301949318, 16.3051294088366, 16.3051288192652, 16.3051284262175, 
    16.3051282296937, 16.3051282296937, 16.3051284262175, 16.3051288192652, 
    16.3051294088366, 16.3051301949318, 16.3051311775506, 16.3051323566929, 
    16.3051337323587, 16.3051353045477, 16.3051370732599, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282, 18.3051282051282, 18.3051282051282, 
    18.3051282051282, 18.3051282051282,
  17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 15.7923165604394, 
    15.7923147917272, 15.7923132195382, 15.7923118438724, 15.79231066473, 
    15.7923096821112, 15.7923088960161, 15.7923083064447, 15.792307913397, 
    15.7923077168732, 15.7923077168732, 15.792307913397, 15.7923083064447, 
    15.7923088960161, 15.7923096821112, 15.79231066473, 15.7923118438724, 
    15.7923132195382, 15.7923147917272, 15.7923165604394, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077,
  17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 15.7923165604394, 
    15.7923147917272, 15.7923132195382, 15.7923118438724, 15.79231066473, 
    15.7923096821112, 15.7923088960161, 15.7923083064447, 15.792307913397, 
    15.7923077168732, 15.7923077168732, 15.792307913397, 15.7923083064447, 
    15.7923088960161, 15.7923096821112, 15.79231066473, 15.7923118438724, 
    15.7923132195382, 15.7923147917272, 15.7923165604394, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077,
  17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 15.7923165604394, 
    15.7923147917272, 15.7923132195382, 15.7923118438724, 15.79231066473, 
    15.7923096821112, 15.7923088960161, 15.7923083064447, 15.792307913397, 
    15.7923077168732, 15.7923077168732, 15.792307913397, 15.7923083064447, 
    15.7923088960161, 15.7923096821112, 15.79231066473, 15.7923118438724, 
    15.7923132195382, 15.7923147917272, 15.7923165604394, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077,
  17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 15.7923165604394, 
    15.7923147917272, 15.7923132195382, 15.7923118438724, 15.79231066473, 
    15.7923096821112, 15.7923088960161, 15.7923083064447, 15.792307913397, 
    15.7923077168732, 15.7923077168732, 15.792307913397, 15.7923083064447, 
    15.7923088960161, 15.7923096821112, 15.79231066473, 15.7923118438724, 
    15.7923132195382, 15.7923147917272, 15.7923165604394, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077, 17.7923076923077, 17.7923076923077, 
    17.7923076923077, 17.7923076923077,
  17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 15.2794960476189, 
    15.2794942789067, 15.2794927067176, 15.2794913310519, 15.2794901519095, 
    15.2794891692907, 15.2794883831956, 15.2794877936241, 15.2794874005765, 
    15.2794872040527, 15.2794872040527, 15.2794874005765, 15.2794877936241, 
    15.2794883831956, 15.2794891692907, 15.2794901519095, 15.2794913310519, 
    15.2794927067176, 15.2794942789067, 15.2794960476189, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872,
  17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 15.2794960476189, 
    15.2794942789067, 15.2794927067176, 15.2794913310519, 15.2794901519095, 
    15.2794891692907, 15.2794883831956, 15.2794877936241, 15.2794874005765, 
    15.2794872040527, 15.2794872040527, 15.2794874005765, 15.2794877936241, 
    15.2794883831956, 15.2794891692907, 15.2794901519095, 15.2794913310519, 
    15.2794927067176, 15.2794942789067, 15.2794960476189, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872,
  17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 15.2794960476189, 
    15.2794942789067, 15.2794927067176, 15.2794913310519, 15.2794901519095, 
    15.2794891692907, 15.2794883831956, 15.2794877936241, 15.2794874005765, 
    15.2794872040527, 15.2794872040527, 15.2794874005765, 15.2794877936241, 
    15.2794883831956, 15.2794891692907, 15.2794901519095, 15.2794913310519, 
    15.2794927067176, 15.2794942789067, 15.2794960476189, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872,
  17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 15.2794960476189, 
    15.2794942789067, 15.2794927067176, 15.2794913310519, 15.2794901519095, 
    15.2794891692907, 15.2794883831956, 15.2794877936241, 15.2794874005765, 
    15.2794872040527, 15.2794872040527, 15.2794874005765, 15.2794877936241, 
    15.2794883831956, 15.2794891692907, 15.2794901519095, 15.2794913310519, 
    15.2794927067176, 15.2794942789067, 15.2794960476189, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872, 17.2794871794872, 17.2794871794872, 
    17.2794871794872, 17.2794871794872,
  16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 14.7666755347984, 
    14.7666737660862, 14.7666721938971, 14.7666708182314, 14.766669639089, 
    14.7666686564702, 14.7666678703751, 14.7666672808036, 14.766666887756, 
    14.7666666912321, 14.7666666912321, 14.766666887756, 14.7666672808036, 
    14.7666678703751, 14.7666686564702, 14.766669639089, 14.7666708182314, 
    14.7666721938971, 14.7666737660862, 14.7666755347984, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667,
  16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 14.7666755347984, 
    14.7666737660862, 14.7666721938971, 14.7666708182314, 14.766669639089, 
    14.7666686564702, 14.7666678703751, 14.7666672808036, 14.766666887756, 
    14.7666666912321, 14.7666666912321, 14.766666887756, 14.7666672808036, 
    14.7666678703751, 14.7666686564702, 14.766669639089, 14.7666708182314, 
    14.7666721938971, 14.7666737660862, 14.7666755347984, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667,
  16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 14.7666755347984, 
    14.7666737660862, 14.7666721938971, 14.7666708182314, 14.766669639089, 
    14.7666686564702, 14.7666678703751, 14.7666672808036, 14.766666887756, 
    14.7666666912321, 14.7666666912321, 14.766666887756, 14.7666672808036, 
    14.7666678703751, 14.7666686564702, 14.766669639089, 14.7666708182314, 
    14.7666721938971, 14.7666737660862, 14.7666755347984, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667,
  16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 14.7666755347984, 
    14.7666737660862, 14.7666721938971, 14.7666708182314, 14.766669639089, 
    14.7666686564702, 14.7666678703751, 14.7666672808036, 14.766666887756, 
    14.7666666912321, 14.7666666912321, 14.766666887756, 14.7666672808036, 
    14.7666678703751, 14.7666686564702, 14.766669639089, 14.7666708182314, 
    14.7666721938971, 14.7666737660862, 14.7666755347984, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667, 16.7666666666667, 16.7666666666667, 
    16.7666666666667, 16.7666666666667,
  16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 14.2538550219779, 
    14.2538532532657, 14.2538516810766, 14.2538503054108, 14.2538491262685, 
    14.2538481436497, 14.2538473575546, 14.2538467679831, 14.2538463749355, 
    14.2538461784116, 14.2538461784116, 14.2538463749355, 14.2538467679831, 
    14.2538473575546, 14.2538481436497, 14.2538491262685, 14.2538503054108, 
    14.2538516810766, 14.2538532532657, 14.2538550219779, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462,
  16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 14.2538550219779, 
    14.2538532532657, 14.2538516810766, 14.2538503054108, 14.2538491262685, 
    14.2538481436497, 14.2538473575546, 14.2538467679831, 14.2538463749355, 
    14.2538461784116, 14.2538461784116, 14.2538463749355, 14.2538467679831, 
    14.2538473575546, 14.2538481436497, 14.2538491262685, 14.2538503054108, 
    14.2538516810766, 14.2538532532657, 14.2538550219779, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462,
  16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 14.2538550219779, 
    14.2538532532657, 14.2538516810766, 14.2538503054108, 14.2538491262685, 
    14.2538481436497, 14.2538473575546, 14.2538467679831, 14.2538463749355, 
    14.2538461784116, 14.2538461784116, 14.2538463749355, 14.2538467679831, 
    14.2538473575546, 14.2538481436497, 14.2538491262685, 14.2538503054108, 
    14.2538516810766, 14.2538532532657, 14.2538550219779, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462,
  16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 14.2538550219779, 
    14.2538532532657, 14.2538516810766, 14.2538503054108, 14.2538491262685, 
    14.2538481436497, 14.2538473575546, 14.2538467679831, 14.2538463749355, 
    14.2538461784116, 14.2538461784116, 14.2538463749355, 14.2538467679831, 
    14.2538473575546, 14.2538481436497, 14.2538491262685, 14.2538503054108, 
    14.2538516810766, 14.2538532532657, 14.2538550219779, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462, 16.2538461538462, 16.2538461538462, 
    16.2538461538462, 16.2538461538462,
  15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 13.7410345091574, 
    13.7410327404452, 13.7410311682561, 13.7410297925903, 13.741028613448, 
    13.7410276308292, 13.741026844734, 13.7410262551626, 13.741025862115, 
    13.7410256655911, 13.7410256655911, 13.741025862115, 13.7410262551626, 
    13.741026844734, 13.7410276308292, 13.741028613448, 13.7410297925903, 
    13.7410311682561, 13.7410327404452, 13.7410345091574, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256,
  15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 13.7410345091574, 
    13.7410327404452, 13.7410311682561, 13.7410297925903, 13.741028613448, 
    13.7410276308292, 13.741026844734, 13.7410262551626, 13.741025862115, 
    13.7410256655911, 13.7410256655911, 13.741025862115, 13.7410262551626, 
    13.741026844734, 13.7410276308292, 13.741028613448, 13.7410297925903, 
    13.7410311682561, 13.7410327404452, 13.7410345091574, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256,
  15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 13.7410345091574, 
    13.7410327404452, 13.7410311682561, 13.7410297925903, 13.741028613448, 
    13.7410276308292, 13.741026844734, 13.7410262551626, 13.741025862115, 
    13.7410256655911, 13.7410256655911, 13.741025862115, 13.7410262551626, 
    13.741026844734, 13.7410276308292, 13.741028613448, 13.7410297925903, 
    13.7410311682561, 13.7410327404452, 13.7410345091574, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256,
  15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 13.7410345091574, 
    13.7410327404452, 13.7410311682561, 13.7410297925903, 13.741028613448, 
    13.7410276308292, 13.741026844734, 13.7410262551626, 13.741025862115, 
    13.7410256655911, 13.7410256655911, 13.741025862115, 13.7410262551626, 
    13.741026844734, 13.7410276308292, 13.741028613448, 13.7410297925903, 
    13.7410311682561, 13.7410327404452, 13.7410345091574, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256, 15.7410256410256, 15.7410256410256, 
    15.7410256410256, 15.7410256410256,
  15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 13.2282139963369, 
    13.2282122276247, 13.2282106554356, 13.2282092797698, 13.2282081006275, 
    13.2282071180087, 13.2282063319135, 13.2282057423421, 13.2282053492944, 
    13.2282051527706, 13.2282051527706, 13.2282053492944, 13.2282057423421, 
    13.2282063319135, 13.2282071180087, 13.2282081006275, 13.2282092797698, 
    13.2282106554356, 13.2282122276247, 13.2282139963369, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051,
  15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 13.2282139963369, 
    13.2282122276247, 13.2282106554356, 13.2282092797698, 13.2282081006275, 
    13.2282071180087, 13.2282063319135, 13.2282057423421, 13.2282053492944, 
    13.2282051527706, 13.2282051527706, 13.2282053492944, 13.2282057423421, 
    13.2282063319135, 13.2282071180087, 13.2282081006275, 13.2282092797698, 
    13.2282106554356, 13.2282122276247, 13.2282139963369, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051,
  15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 13.2282139963369, 
    13.2282122276247, 13.2282106554356, 13.2282092797698, 13.2282081006275, 
    13.2282071180087, 13.2282063319135, 13.2282057423421, 13.2282053492944, 
    13.2282051527706, 13.2282051527706, 13.2282053492944, 13.2282057423421, 
    13.2282063319135, 13.2282071180087, 13.2282081006275, 13.2282092797698, 
    13.2282106554356, 13.2282122276247, 13.2282139963369, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051,
  15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 13.2282139963369, 
    13.2282122276247, 13.2282106554356, 13.2282092797698, 13.2282081006275, 
    13.2282071180087, 13.2282063319135, 13.2282057423421, 13.2282053492944, 
    13.2282051527706, 13.2282051527706, 13.2282053492944, 13.2282057423421, 
    13.2282063319135, 13.2282071180087, 13.2282081006275, 13.2282092797698, 
    13.2282106554356, 13.2282122276247, 13.2282139963369, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051, 15.2282051282051, 15.2282051282051, 
    15.2282051282051, 15.2282051282051,
  14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 12.7153934835164, 
    12.7153917148041, 12.7153901426151, 12.7153887669493, 12.715387587807, 
    12.7153866051882, 12.715385819093, 12.7153852295216, 12.7153848364739, 
    12.7153846399501, 12.7153846399501, 12.7153848364739, 12.7153852295216, 
    12.715385819093, 12.7153866051882, 12.715387587807, 12.7153887669493, 
    12.7153901426151, 12.7153917148041, 12.7153934835164, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846,
  14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 12.7153934835164, 
    12.7153917148041, 12.7153901426151, 12.7153887669493, 12.715387587807, 
    12.7153866051882, 12.715385819093, 12.7153852295216, 12.7153848364739, 
    12.7153846399501, 12.7153846399501, 12.7153848364739, 12.7153852295216, 
    12.715385819093, 12.7153866051882, 12.715387587807, 12.7153887669493, 
    12.7153901426151, 12.7153917148041, 12.7153934835164, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846,
  14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 12.7153934835164, 
    12.7153917148041, 12.7153901426151, 12.7153887669493, 12.715387587807, 
    12.7153866051882, 12.715385819093, 12.7153852295216, 12.7153848364739, 
    12.7153846399501, 12.7153846399501, 12.7153848364739, 12.7153852295216, 
    12.715385819093, 12.7153866051882, 12.715387587807, 12.7153887669493, 
    12.7153901426151, 12.7153917148041, 12.7153934835164, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846,
  14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 12.7153934835164, 
    12.7153917148041, 12.7153901426151, 12.7153887669493, 12.715387587807, 
    12.7153866051882, 12.715385819093, 12.7153852295216, 12.7153848364739, 
    12.7153846399501, 12.7153846399501, 12.7153848364739, 12.7153852295216, 
    12.715385819093, 12.7153866051882, 12.715387587807, 12.7153887669493, 
    12.7153901426151, 12.7153917148041, 12.7153934835164, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846, 14.7153846153846, 14.7153846153846, 
    14.7153846153846, 14.7153846153846,
  14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 12.2025729706958, 
    12.2025712019836, 12.2025696297946, 12.2025682541288, 12.2025670749865, 
    12.2025660923677, 12.2025653062725, 12.2025647167011, 12.2025643236534, 
    12.2025641271296, 12.2025641271296, 12.2025643236534, 12.2025647167011, 
    12.2025653062725, 12.2025660923677, 12.2025670749865, 12.2025682541288, 
    12.2025696297946, 12.2025712019836, 12.2025729706958, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641,
  14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 12.2025729706958, 
    12.2025712019836, 12.2025696297946, 12.2025682541288, 12.2025670749865, 
    12.2025660923677, 12.2025653062725, 12.2025647167011, 12.2025643236534, 
    12.2025641271296, 12.2025641271296, 12.2025643236534, 12.2025647167011, 
    12.2025653062725, 12.2025660923677, 12.2025670749865, 12.2025682541288, 
    12.2025696297946, 12.2025712019836, 12.2025729706958, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641,
  14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 12.2025729706958, 
    12.2025712019836, 12.2025696297946, 12.2025682541288, 12.2025670749865, 
    12.2025660923677, 12.2025653062725, 12.2025647167011, 12.2025643236534, 
    12.2025641271296, 12.2025641271296, 12.2025643236534, 12.2025647167011, 
    12.2025653062725, 12.2025660923677, 12.2025670749865, 12.2025682541288, 
    12.2025696297946, 12.2025712019836, 12.2025729706958, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641,
  14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 12.2025729706958, 
    12.2025712019836, 12.2025696297946, 12.2025682541288, 12.2025670749865, 
    12.2025660923677, 12.2025653062725, 12.2025647167011, 12.2025643236534, 
    12.2025641271296, 12.2025641271296, 12.2025643236534, 12.2025647167011, 
    12.2025653062725, 12.2025660923677, 12.2025670749865, 12.2025682541288, 
    12.2025696297946, 12.2025712019836, 12.2025729706958, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641, 14.2025641025641, 14.2025641025641, 
    14.2025641025641, 14.2025641025641,
  13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 11.6897524578753, 
    11.6897506891631, 11.6897491169741, 11.6897477413083, 11.6897465621659, 
    11.6897455795471, 11.689744793452, 11.6897442038806, 11.6897438108329, 
    11.6897436143091, 11.6897436143091, 11.6897438108329, 11.6897442038806, 
    11.689744793452, 11.6897455795471, 11.6897465621659, 11.6897477413083, 
    11.6897491169741, 11.6897506891631, 11.6897524578753, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436,
  13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 11.6897524578753, 
    11.6897506891631, 11.6897491169741, 11.6897477413083, 11.6897465621659, 
    11.6897455795471, 11.689744793452, 11.6897442038806, 11.6897438108329, 
    11.6897436143091, 11.6897436143091, 11.6897438108329, 11.6897442038806, 
    11.689744793452, 11.6897455795471, 11.6897465621659, 11.6897477413083, 
    11.6897491169741, 11.6897506891631, 11.6897524578753, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436,
  13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 11.6897524578753, 
    11.6897506891631, 11.6897491169741, 11.6897477413083, 11.6897465621659, 
    11.6897455795471, 11.689744793452, 11.6897442038806, 11.6897438108329, 
    11.6897436143091, 11.6897436143091, 11.6897438108329, 11.6897442038806, 
    11.689744793452, 11.6897455795471, 11.6897465621659, 11.6897477413083, 
    11.6897491169741, 11.6897506891631, 11.6897524578753, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436,
  13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 11.6897524578753, 
    11.6897506891631, 11.6897491169741, 11.6897477413083, 11.6897465621659, 
    11.6897455795471, 11.689744793452, 11.6897442038806, 11.6897438108329, 
    11.6897436143091, 11.6897436143091, 11.6897438108329, 11.6897442038806, 
    11.689744793452, 11.6897455795471, 11.6897465621659, 11.6897477413083, 
    11.6897491169741, 11.6897506891631, 11.6897524578753, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436, 13.6897435897436, 13.6897435897436, 
    13.6897435897436, 13.6897435897436,
  13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 11.1769319450548, 
    11.1769301763426, 11.1769286041535, 11.1769272284878, 11.1769260493454, 
    11.1769250667266, 11.1769242806315, 11.17692369106, 11.1769232980124, 
    11.1769231014886, 11.1769231014886, 11.1769232980124, 11.17692369106, 
    11.1769242806315, 11.1769250667266, 11.1769260493454, 11.1769272284878, 
    11.1769286041535, 11.1769301763426, 11.1769319450548, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231,
  13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 11.1769319450548, 
    11.1769301763426, 11.1769286041535, 11.1769272284878, 11.1769260493454, 
    11.1769250667266, 11.1769242806315, 11.17692369106, 11.1769232980124, 
    11.1769231014886, 11.1769231014886, 11.1769232980124, 11.17692369106, 
    11.1769242806315, 11.1769250667266, 11.1769260493454, 11.1769272284878, 
    11.1769286041535, 11.1769301763426, 11.1769319450548, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231,
  13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 11.1769319450548, 
    11.1769301763426, 11.1769286041535, 11.1769272284878, 11.1769260493454, 
    11.1769250667266, 11.1769242806315, 11.17692369106, 11.1769232980124, 
    11.1769231014886, 11.1769231014886, 11.1769232980124, 11.17692369106, 
    11.1769242806315, 11.1769250667266, 11.1769260493454, 11.1769272284878, 
    11.1769286041535, 11.1769301763426, 11.1769319450548, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231,
  13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 11.1769319450548, 
    11.1769301763426, 11.1769286041535, 11.1769272284878, 11.1769260493454, 
    11.1769250667266, 11.1769242806315, 11.17692369106, 11.1769232980124, 
    11.1769231014886, 11.1769231014886, 11.1769232980124, 11.17692369106, 
    11.1769242806315, 11.1769250667266, 11.1769260493454, 11.1769272284878, 
    11.1769286041535, 11.1769301763426, 11.1769319450548, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231, 13.1769230769231, 13.1769230769231, 
    13.1769230769231, 13.1769230769231,
  12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 10.6641114322343, 
    10.6641096635221, 10.664108091333, 10.6641067156673, 10.6641055365249, 
    10.6641045539061, 10.664103767811, 10.6641031782395, 10.6641027851919, 
    10.664102588668, 10.664102588668, 10.6641027851919, 10.6641031782395, 
    10.664103767811, 10.6641045539061, 10.6641055365249, 10.6641067156673, 
    10.664108091333, 10.6641096635221, 10.6641114322343, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026,
  12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 10.6641114322343, 
    10.6641096635221, 10.664108091333, 10.6641067156673, 10.6641055365249, 
    10.6641045539061, 10.664103767811, 10.6641031782395, 10.6641027851919, 
    10.664102588668, 10.664102588668, 10.6641027851919, 10.6641031782395, 
    10.664103767811, 10.6641045539061, 10.6641055365249, 10.6641067156673, 
    10.664108091333, 10.6641096635221, 10.6641114322343, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026,
  12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 10.6641114322343, 
    10.6641096635221, 10.664108091333, 10.6641067156673, 10.6641055365249, 
    10.6641045539061, 10.664103767811, 10.6641031782395, 10.6641027851919, 
    10.664102588668, 10.664102588668, 10.6641027851919, 10.6641031782395, 
    10.664103767811, 10.6641045539061, 10.6641055365249, 10.6641067156673, 
    10.664108091333, 10.6641096635221, 10.6641114322343, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026,
  12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 10.6641114322343, 
    10.6641096635221, 10.664108091333, 10.6641067156673, 10.6641055365249, 
    10.6641045539061, 10.664103767811, 10.6641031782395, 10.6641027851919, 
    10.664102588668, 10.664102588668, 10.6641027851919, 10.6641031782395, 
    10.664103767811, 10.6641045539061, 10.6641055365249, 10.6641067156673, 
    10.664108091333, 10.6641096635221, 10.6641114322343, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026, 12.6641025641026, 12.6641025641026, 
    12.6641025641026, 12.6641025641026,
  12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 10.1512909194138, 
    10.1512891507016, 10.1512875785125, 10.1512862028467, 10.1512850237044, 
    10.1512840410856, 10.1512832549905, 10.151282665419, 10.1512822723714, 
    10.1512820758475, 10.1512820758475, 10.1512822723714, 10.151282665419, 
    10.1512832549905, 10.1512840410856, 10.1512850237044, 10.1512862028467, 
    10.1512875785125, 10.1512891507016, 10.1512909194138, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821,
  12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 10.1512909194138, 
    10.1512891507016, 10.1512875785125, 10.1512862028467, 10.1512850237044, 
    10.1512840410856, 10.1512832549905, 10.151282665419, 10.1512822723714, 
    10.1512820758475, 10.1512820758475, 10.1512822723714, 10.151282665419, 
    10.1512832549905, 10.1512840410856, 10.1512850237044, 10.1512862028467, 
    10.1512875785125, 10.1512891507016, 10.1512909194138, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821,
  12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 10.1512909194138, 
    10.1512891507016, 10.1512875785125, 10.1512862028467, 10.1512850237044, 
    10.1512840410856, 10.1512832549905, 10.151282665419, 10.1512822723714, 
    10.1512820758475, 10.1512820758475, 10.1512822723714, 10.151282665419, 
    10.1512832549905, 10.1512840410856, 10.1512850237044, 10.1512862028467, 
    10.1512875785125, 10.1512891507016, 10.1512909194138, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821,
  12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 10.1512909194138, 
    10.1512891507016, 10.1512875785125, 10.1512862028467, 10.1512850237044, 
    10.1512840410856, 10.1512832549905, 10.151282665419, 10.1512822723714, 
    10.1512820758475, 10.1512820758475, 10.1512822723714, 10.151282665419, 
    10.1512832549905, 10.1512840410856, 10.1512850237044, 10.1512862028467, 
    10.1512875785125, 10.1512891507016, 10.1512909194138, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821, 12.1512820512821, 12.1512820512821, 
    12.1512820512821, 12.1512820512821,
  11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 9.63847040659328, 
    9.63846863788107, 9.638467065692, 9.63846569002623, 9.63846451088389, 
    9.63846352826509, 9.63846274216994, 9.63846215259851, 9.63846175955085, 
    9.63846156302702, 9.63846156302702, 9.63846175955085, 9.63846215259851, 
    9.63846274216994, 9.63846352826509, 9.63846451088389, 9.63846569002623, 
    9.638467065692, 9.63846863788107, 9.63847040659328, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615,
  11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 9.63847040659328, 
    9.63846863788107, 9.638467065692, 9.63846569002623, 9.63846451088389, 
    9.63846352826509, 9.63846274216994, 9.63846215259851, 9.63846175955085, 
    9.63846156302702, 9.63846156302702, 9.63846175955085, 9.63846215259851, 
    9.63846274216994, 9.63846352826509, 9.63846451088389, 9.63846569002623, 
    9.638467065692, 9.63846863788107, 9.63847040659328, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615,
  11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 9.63847040659328, 
    9.63846863788107, 9.638467065692, 9.63846569002623, 9.63846451088389, 
    9.63846352826509, 9.63846274216994, 9.63846215259851, 9.63846175955085, 
    9.63846156302702, 9.63846156302702, 9.63846175955085, 9.63846215259851, 
    9.63846274216994, 9.63846352826509, 9.63846451088389, 9.63846569002623, 
    9.638467065692, 9.63846863788107, 9.63847040659328, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615,
  11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 9.63847040659328, 
    9.63846863788107, 9.638467065692, 9.63846569002623, 9.63846451088389, 
    9.63846352826509, 9.63846274216994, 9.63846215259851, 9.63846175955085, 
    9.63846156302702, 9.63846156302702, 9.63846175955085, 9.63846215259851, 
    9.63846274216994, 9.63846352826509, 9.63846451088389, 9.63846569002623, 
    9.638467065692, 9.63846863788107, 9.63847040659328, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615, 11.6384615384615, 11.6384615384615, 
    11.6384615384615, 11.6384615384615,
  11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 9.12564989377277, 
    9.12564812506056, 9.12564655287149, 9.12564517720572, 9.12564399806337, 
    9.12564301544458, 9.12564222934943, 9.125641639778, 9.12564124673034, 
    9.12564105020651, 9.12564105020651, 9.12564124673034, 9.125641639778, 
    9.12564222934943, 9.12564301544458, 9.12564399806337, 9.12564517720572, 
    9.12564655287149, 9.12564812506056, 9.12564989377277, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641,
  11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 9.12564989377277, 
    9.12564812506056, 9.12564655287149, 9.12564517720572, 9.12564399806337, 
    9.12564301544458, 9.12564222934943, 9.125641639778, 9.12564124673034, 
    9.12564105020651, 9.12564105020651, 9.12564124673034, 9.125641639778, 
    9.12564222934943, 9.12564301544458, 9.12564399806337, 9.12564517720572, 
    9.12564655287149, 9.12564812506056, 9.12564989377277, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641,
  11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 9.12564989377277, 
    9.12564812506056, 9.12564655287149, 9.12564517720572, 9.12564399806337, 
    9.12564301544458, 9.12564222934943, 9.125641639778, 9.12564124673034, 
    9.12564105020651, 9.12564105020651, 9.12564124673034, 9.125641639778, 
    9.12564222934943, 9.12564301544458, 9.12564399806337, 9.12564517720572, 
    9.12564655287149, 9.12564812506056, 9.12564989377277, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641,
  11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 9.12564989377277, 
    9.12564812506056, 9.12564655287149, 9.12564517720572, 9.12564399806337, 
    9.12564301544458, 9.12564222934943, 9.125641639778, 9.12564124673034, 
    9.12564105020651, 9.12564105020651, 9.12564124673034, 9.125641639778, 
    9.12564222934943, 9.12564301544458, 9.12564399806337, 9.12564517720572, 
    9.12564655287149, 9.12564812506056, 9.12564989377277, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641, 11.125641025641, 11.125641025641, 
    11.125641025641, 11.125641025641,
  10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 8.61282938095225, 
    8.61282761224004, 8.61282604005098, 8.6128246643852, 8.61282348524286, 
    8.61282250262407, 8.61282171652891, 8.61282112695748, 8.61282073390983, 
    8.61282053738599, 8.61282053738599, 8.61282073390983, 8.61282112695748, 
    8.61282171652891, 8.61282250262407, 8.61282348524286, 8.6128246643852, 
    8.61282604005098, 8.61282761224004, 8.61282938095225, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205,
  10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 8.61282938095225, 
    8.61282761224004, 8.61282604005098, 8.6128246643852, 8.61282348524286, 
    8.61282250262407, 8.61282171652891, 8.61282112695748, 8.61282073390983, 
    8.61282053738599, 8.61282053738599, 8.61282073390983, 8.61282112695748, 
    8.61282171652891, 8.61282250262407, 8.61282348524286, 8.6128246643852, 
    8.61282604005098, 8.61282761224004, 8.61282938095225, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205,
  10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 8.61282938095225, 
    8.61282761224004, 8.61282604005098, 8.6128246643852, 8.61282348524286, 
    8.61282250262407, 8.61282171652891, 8.61282112695748, 8.61282073390983, 
    8.61282053738599, 8.61282053738599, 8.61282073390983, 8.61282112695748, 
    8.61282171652891, 8.61282250262407, 8.61282348524286, 8.6128246643852, 
    8.61282604005098, 8.61282761224004, 8.61282938095225, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205,
  10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 8.61282938095225, 
    8.61282761224004, 8.61282604005098, 8.6128246643852, 8.61282348524286, 
    8.61282250262407, 8.61282171652891, 8.61282112695748, 8.61282073390983, 
    8.61282053738599, 8.61282053738599, 8.61282073390983, 8.61282112695748, 
    8.61282171652891, 8.61282250262407, 8.61282348524286, 8.6128246643852, 
    8.61282604005098, 8.61282761224004, 8.61282938095225, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205, 10.6128205128205, 10.6128205128205, 
    10.6128205128205, 10.6128205128205,
  10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 8.10000886813174, 8.10000709941953, 8.10000552723046, 
    8.10000415156469, 8.10000297242235, 8.10000198980355, 8.1000012037084, 
    8.10000061413697, 8.10000022108932, 8.10000002456548, 8.10000002456548, 
    8.10000022108932, 8.10000061413697, 8.1000012037084, 8.10000198980355, 
    8.10000297242235, 8.10000415156469, 8.10000552723046, 8.10000709941953, 
    8.10000886813174, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1,
  10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 8.10000886813174, 8.10000709941953, 8.10000552723046, 
    8.10000415156469, 8.10000297242235, 8.10000198980355, 8.1000012037084, 
    8.10000061413697, 8.10000022108932, 8.10000002456548, 8.10000002456548, 
    8.10000022108932, 8.10000061413697, 8.1000012037084, 8.10000198980355, 
    8.10000297242235, 8.10000415156469, 8.10000552723046, 8.10000709941953, 
    8.10000886813174, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1,
  10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 8.10000886813174, 8.10000709941953, 8.10000552723046, 
    8.10000415156469, 8.10000297242235, 8.10000198980355, 8.1000012037084, 
    8.10000061413697, 8.10000022108932, 8.10000002456548, 8.10000002456548, 
    8.10000022108932, 8.10000061413697, 8.1000012037084, 8.10000198980355, 
    8.10000297242235, 8.10000415156469, 8.10000552723046, 8.10000709941953, 
    8.10000886813174, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1,
  10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 8.10000886813174, 8.10000709941953, 8.10000552723046, 
    8.10000415156469, 8.10000297242235, 8.10000198980355, 8.1000012037084, 
    8.10000061413697, 8.10000022108932, 8.10000002456548, 8.10000002456548, 
    8.10000022108932, 8.10000061413697, 8.1000012037084, 8.10000198980355, 
    8.10000297242235, 8.10000415156469, 8.10000552723046, 8.10000709941953, 
    8.10000886813174, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 10.1, 
    10.1, 10.1, 10.1, 10.1, 10.1, 10.1 ;

 salt =
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35 ;
}
